module AN2(a, b, z);

input	a, b;
output	z;

and #1 g1(z, a, b);

endmodule
