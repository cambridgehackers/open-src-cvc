module	OR2(a, b, z);

input	a, b;
output	z;

or #1 g1(z, a, b);

endmodule
