// DA Solutions Ltd., Testbench to drive DA Solutions provided
// Multiplier circuit
// Creeated 1-Sep-94, D. J. Wharton
// Circuit also available in VHDL
// Library used LCA100k CMOS
 
`timescale 1ns / 10 ps
module testbench;

reg	[0:112]	patternsin[0:3095];
reg	[0:112] inbuf1, inbuf2;
reg	[8:63]	patternsout[0:1547];
reg	[8:63]	outbuf;
reg	[0:63]	errorbit;

reg	[8:63]	oper1, oper2;
reg		do_mult;

wire	[8:63]	product;

initial
begin
//	$readmemb ("/home/vecircs/DAS/mult/ref_in", patternsin);
	$readmemb ("ref_in", patternsin);
//	$readmemb ("/home/vecircs/DAS/mult/ref_out", patternsout);
	$readmemb ("ref_out", patternsout);
	do_mult = 1;
	begin : multpattloop
	integer i;
	for (i=0; i < 3096; i = i + 2)
	begin
	   #5	do_mult = 0;
	   #95	inbuf1 = patternsin[i];
		inbuf2 = patternsin[i+1];
		oper1 = inbuf1;
		oper2 = inbuf2;
		outbuf = patternsout[i/2];
	   #5	do_mult =1;
	   #395	errorbit = product ^ outbuf;
		if (errorbit != 0)
			begin
			$display ($time,,,,"Output miscompare");
			$display ($time,,,,"error register =",,errorbit,,,,"prod",,product,,,,"buf",,outbuf,,,,"loopcount",,i);
			end
	end
	end
end

mult_56		component1 (oper1, oper2, product, do_mult);

endmodule

// End of testbench


// Author	D. J. Wharton, DA Solutions Ltd
// Date		1-Sep-94
// Version 	1.0
// File		mult_56_gate.v
// Gate level version of 56 bit floating point multiplier

module	mult_56 (oper1[8:63], oper2[8:63], product[8:63], do_mult);

input	[8:63]	oper1, oper2;
output	[8:63]	product;
input		do_mult;
wire	[8:63]	gen, tr,carry; //, g63;
wire	[0:7]	ggen, gtran, gcarry;
wire	[8:63]	nop;

wire	[8:63]	g63, g62, g61, g60, g59, g58, g57, g56;
wire	[8:63]	g55, g54, g53, g52, g51, g50, g49, g48;
wire	[8:63]	g47, g46, g45, g44, g43, g42, g41, g40;
wire	[8:63]	g39, g38, g37, g36, g35, g34, g33, g32;
wire	[8:63]	g31, g30, g29, g28, g27, g26, g25, g24;
wire	[8:63]	g23, g22, g21, g20, g19, g18, g17, g16;
wire	[8:63]	g15, g14, g13, g12, g11, g10, g9, g8;

wire    [8:63]  pc63, pc62, pc61, pc60, pc59, pc58, pc57, pc56;
wire    [8:63]  pc55, pc54, pc53, pc52, pc51, pc50, pc49, pc48;
wire    [8:63]  pc47, pc46, pc45, pc44, pc43, pc42, pc41, pc40;
wire    [8:63]  pc39, pc38, pc37, pc36, pc35, pc34, pc33, pc32;
wire    [8:63]  pc31, pc30, pc29, pc28, pc27, pc26, pc25, pc24;
wire    [8:63]  pc23, pc22, pc21, pc20, pc19, pc18, pc17, pc16;
wire    [8:63]  pc15, pc14, pc13, pc12, pc11, pc10, pc9, pc8;

wire    [8:63]  ps63, ps62, ps61, ps60, ps59, ps58, ps57, ps56;
wire    [8:63]  ps55, ps54, ps53, ps52, ps51, ps50, ps49, ps48;
wire    [8:63]  ps47, ps46, ps45, ps44, ps43, ps42, ps41, ps40;
wire    [8:63]  ps39, ps38, ps37, ps36, ps35, ps34, ps33, ps32;
wire    [8:63]  ps31, ps30, ps29, ps28, ps27, ps26, ps25, ps24;
wire    [8:63]  ps23, ps22, ps21, ps20, ps19, ps18, ps17, ps16;
wire    [8:63]  ps15, ps14, ps13, ps12, ps11, ps10, ps9, ps8;


`define	zero 1'b0

carry_block GCB1(gen[8:15], tr[8:15], carry[8:15], gcarry[0], ggen[0], gtran[0]);
carry_block GCB2(gen[16:23], tr[16:23], carry[16:23], gcarry[1], ggen[1], gtran[1]);
carry_block GCB3(gen[24:31], tr[24:31], carry[24:31], gcarry[2], ggen[2], gtran[2]);
carry_block GCB4(gen[32:39], tr[32:39], carry[32:39], gcarry[3], ggen[3], gtran[3]);
carry_block GCB5(gen[40:47], tr[40:47], carry[40:47], gcarry[4], ggen[4], gtran[4]);
carry_block GCB6(gen[48:55], tr[48:55], carry[48:55], gcarry[5], ggen[5], gtran[5]);
carry_block GCB7(gen[56:63], tr[56:63], carry[56:63], `zero, ggen[6], gtran[6]);
carry_block GGCB(ggen[0:7], gtran[0:7], gcarry[0:7], `zero, ggg, ggt);
BUF8A GB1(`zero, gen[63]);
BUF8A GB2(`zero, tr[63]);
BUF8A GB3(`zero, ggen[7]);
BUF8A GB4(`zero, gtran[7]);
AN2 GA63_8(oper2[8], oper1[63], g63[8]);
AN2 GA63_9(oper2[9], oper1[63], g63[9]);
AN2 GA63_10(oper2[10], oper1[63], g63[10]);
AN2 GA63_11(oper2[11], oper1[63], g63[11]);
AN2 GA63_12(oper2[12], oper1[63], g63[12]);
AN2 GA63_13(oper2[13], oper1[63], g63[13]);
AN2 GA63_14(oper2[14], oper1[63], g63[14]);
AN2 GA63_15(oper2[15], oper1[63], g63[15]);
AN2 GA63_16(oper2[16], oper1[63], g63[16]);
AN2 GA63_17(oper2[17], oper1[63], g63[17]);
AN2 GA63_18(oper2[18], oper1[63], g63[18]);
AN2 GA63_19(oper2[19], oper1[63], g63[19]);
AN2 GA63_20(oper2[20], oper1[63], g63[20]);
AN2 GA63_21(oper2[21], oper1[63], g63[21]);
AN2 GA63_22(oper2[22], oper1[63], g63[22]);
AN2 GA63_23(oper2[23], oper1[63], g63[23]);
AN2 GA63_24(oper2[24], oper1[63], g63[24]);
AN2 GA63_25(oper2[25], oper1[63], g63[25]);
AN2 GA63_26(oper2[26], oper1[63], g63[26]);
AN2 GA63_27(oper2[27], oper1[63], g63[27]);
AN2 GA63_28(oper2[28], oper1[63], g63[28]);
AN2 GA63_29(oper2[29], oper1[63], g63[29]);
AN2 GA63_30(oper2[30], oper1[63], g63[30]);
AN2 GA63_31(oper2[31], oper1[63], g63[31]);
AN2 GA63_32(oper2[32], oper1[63], g63[32]);
AN2 GA63_33(oper2[33], oper1[63], g63[33]);
AN2 GA63_34(oper2[34], oper1[63], g63[34]);
AN2 GA63_35(oper2[35], oper1[63], g63[35]);
AN2 GA63_36(oper2[36], oper1[63], g63[36]);
AN2 GA63_37(oper2[37], oper1[63], g63[37]);
AN2 GA63_38(oper2[38], oper1[63], g63[38]);
AN2 GA63_39(oper2[39], oper1[63], g63[39]);
AN2 GA63_40(oper2[40], oper1[63], g63[40]);
AN2 GA63_41(oper2[41], oper1[63], g63[41]);
AN2 GA63_42(oper2[42], oper1[63], g63[42]);
AN2 GA63_43(oper2[43], oper1[63], g63[43]);
AN2 GA63_44(oper2[44], oper1[63], g63[44]);
AN2 GA63_45(oper2[45], oper1[63], g63[45]);
AN2 GA63_46(oper2[46], oper1[63], g63[46]);
AN2 GA63_47(oper2[47], oper1[63], g63[47]);
AN2 GA63_48(oper2[48], oper1[63], g63[48]);
AN2 GA63_49(oper2[49], oper1[63], g63[49]);
AN2 GA63_50(oper2[50], oper1[63], g63[50]);
AN2 GA63_51(oper2[51], oper1[63], g63[51]);
AN2 GA63_52(oper2[52], oper1[63], g63[52]);
AN2 GA63_53(oper2[53], oper1[63], g63[53]);
AN2 GA63_54(oper2[54], oper1[63], g63[54]);
AN2 GA63_55(oper2[55], oper1[63], g63[55]);
AN2 GA63_56(oper2[56], oper1[63], g63[56]);
AN2 GA63_57(oper2[57], oper1[63], g63[57]);
AN2 GA63_58(oper2[58], oper1[63], g63[58]);
AN2 GA63_59(oper2[59], oper1[63], g63[59]);
AN2 GA63_60(oper2[60], oper1[63], g63[60]);
AN2 GA63_61(oper2[61], oper1[63], g63[61]);
AN2 GA63_62(oper2[62], oper1[63], g63[62]);
AN2 GA63_63(oper2[63], oper1[63], g63[63]);
AN2 GA62_8(oper2[8], oper1[62], g62[8]);
AN2 GA62_9(oper2[9], oper1[62], g62[9]);
AN2 GA62_10(oper2[10], oper1[62], g62[10]);
AN2 GA62_11(oper2[11], oper1[62], g62[11]);
AN2 GA62_12(oper2[12], oper1[62], g62[12]);
AN2 GA62_13(oper2[13], oper1[62], g62[13]);
AN2 GA62_14(oper2[14], oper1[62], g62[14]);
AN2 GA62_15(oper2[15], oper1[62], g62[15]);
AN2 GA62_16(oper2[16], oper1[62], g62[16]);
AN2 GA62_17(oper2[17], oper1[62], g62[17]);
AN2 GA62_18(oper2[18], oper1[62], g62[18]);
AN2 GA62_19(oper2[19], oper1[62], g62[19]);
AN2 GA62_20(oper2[20], oper1[62], g62[20]);
AN2 GA62_21(oper2[21], oper1[62], g62[21]);
AN2 GA62_22(oper2[22], oper1[62], g62[22]);
AN2 GA62_23(oper2[23], oper1[62], g62[23]);
AN2 GA62_24(oper2[24], oper1[62], g62[24]);
AN2 GA62_25(oper2[25], oper1[62], g62[25]);
AN2 GA62_26(oper2[26], oper1[62], g62[26]);
AN2 GA62_27(oper2[27], oper1[62], g62[27]);
AN2 GA62_28(oper2[28], oper1[62], g62[28]);
AN2 GA62_29(oper2[29], oper1[62], g62[29]);
AN2 GA62_30(oper2[30], oper1[62], g62[30]);
AN2 GA62_31(oper2[31], oper1[62], g62[31]);
AN2 GA62_32(oper2[32], oper1[62], g62[32]);
AN2 GA62_33(oper2[33], oper1[62], g62[33]);
AN2 GA62_34(oper2[34], oper1[62], g62[34]);
AN2 GA62_35(oper2[35], oper1[62], g62[35]);
AN2 GA62_36(oper2[36], oper1[62], g62[36]);
AN2 GA62_37(oper2[37], oper1[62], g62[37]);
AN2 GA62_38(oper2[38], oper1[62], g62[38]);
AN2 GA62_39(oper2[39], oper1[62], g62[39]);
AN2 GA62_40(oper2[40], oper1[62], g62[40]);
AN2 GA62_41(oper2[41], oper1[62], g62[41]);
AN2 GA62_42(oper2[42], oper1[62], g62[42]);
AN2 GA62_43(oper2[43], oper1[62], g62[43]);
AN2 GA62_44(oper2[44], oper1[62], g62[44]);
AN2 GA62_45(oper2[45], oper1[62], g62[45]);
AN2 GA62_46(oper2[46], oper1[62], g62[46]);
AN2 GA62_47(oper2[47], oper1[62], g62[47]);
AN2 GA62_48(oper2[48], oper1[62], g62[48]);
AN2 GA62_49(oper2[49], oper1[62], g62[49]);
AN2 GA62_50(oper2[50], oper1[62], g62[50]);
AN2 GA62_51(oper2[51], oper1[62], g62[51]);
AN2 GA62_52(oper2[52], oper1[62], g62[52]);
AN2 GA62_53(oper2[53], oper1[62], g62[53]);
AN2 GA62_54(oper2[54], oper1[62], g62[54]);
AN2 GA62_55(oper2[55], oper1[62], g62[55]);
AN2 GA62_56(oper2[56], oper1[62], g62[56]);
AN2 GA62_57(oper2[57], oper1[62], g62[57]);
AN2 GA62_58(oper2[58], oper1[62], g62[58]);
AN2 GA62_59(oper2[59], oper1[62], g62[59]);
AN2 GA62_60(oper2[60], oper1[62], g62[60]);
AN2 GA62_61(oper2[61], oper1[62], g62[61]);
AN2 GA62_62(oper2[62], oper1[62], g62[62]);
AN2 GA62_63(oper2[63], oper1[62], g62[63]);
AN2 GA61_8(oper2[8], oper1[61], g61[8]);
AN2 GA61_9(oper2[9], oper1[61], g61[9]);
AN2 GA61_10(oper2[10], oper1[61], g61[10]);
AN2 GA61_11(oper2[11], oper1[61], g61[11]);
AN2 GA61_12(oper2[12], oper1[61], g61[12]);
AN2 GA61_13(oper2[13], oper1[61], g61[13]);
AN2 GA61_14(oper2[14], oper1[61], g61[14]);
AN2 GA61_15(oper2[15], oper1[61], g61[15]);
AN2 GA61_16(oper2[16], oper1[61], g61[16]);
AN2 GA61_17(oper2[17], oper1[61], g61[17]);
AN2 GA61_18(oper2[18], oper1[61], g61[18]);
AN2 GA61_19(oper2[19], oper1[61], g61[19]);
AN2 GA61_20(oper2[20], oper1[61], g61[20]);
AN2 GA61_21(oper2[21], oper1[61], g61[21]);
AN2 GA61_22(oper2[22], oper1[61], g61[22]);
AN2 GA61_23(oper2[23], oper1[61], g61[23]);
AN2 GA61_24(oper2[24], oper1[61], g61[24]);
AN2 GA61_25(oper2[25], oper1[61], g61[25]);
AN2 GA61_26(oper2[26], oper1[61], g61[26]);
AN2 GA61_27(oper2[27], oper1[61], g61[27]);
AN2 GA61_28(oper2[28], oper1[61], g61[28]);
AN2 GA61_29(oper2[29], oper1[61], g61[29]);
AN2 GA61_30(oper2[30], oper1[61], g61[30]);
AN2 GA61_31(oper2[31], oper1[61], g61[31]);
AN2 GA61_32(oper2[32], oper1[61], g61[32]);
AN2 GA61_33(oper2[33], oper1[61], g61[33]);
AN2 GA61_34(oper2[34], oper1[61], g61[34]);
AN2 GA61_35(oper2[35], oper1[61], g61[35]);
AN2 GA61_36(oper2[36], oper1[61], g61[36]);
AN2 GA61_37(oper2[37], oper1[61], g61[37]);
AN2 GA61_38(oper2[38], oper1[61], g61[38]);
AN2 GA61_39(oper2[39], oper1[61], g61[39]);
AN2 GA61_40(oper2[40], oper1[61], g61[40]);
AN2 GA61_41(oper2[41], oper1[61], g61[41]);
AN2 GA61_42(oper2[42], oper1[61], g61[42]);
AN2 GA61_43(oper2[43], oper1[61], g61[43]);
AN2 GA61_44(oper2[44], oper1[61], g61[44]);
AN2 GA61_45(oper2[45], oper1[61], g61[45]);
AN2 GA61_46(oper2[46], oper1[61], g61[46]);
AN2 GA61_47(oper2[47], oper1[61], g61[47]);
AN2 GA61_48(oper2[48], oper1[61], g61[48]);
AN2 GA61_49(oper2[49], oper1[61], g61[49]);
AN2 GA61_50(oper2[50], oper1[61], g61[50]);
AN2 GA61_51(oper2[51], oper1[61], g61[51]);
AN2 GA61_52(oper2[52], oper1[61], g61[52]);
AN2 GA61_53(oper2[53], oper1[61], g61[53]);
AN2 GA61_54(oper2[54], oper1[61], g61[54]);
AN2 GA61_55(oper2[55], oper1[61], g61[55]);
AN2 GA61_56(oper2[56], oper1[61], g61[56]);
AN2 GA61_57(oper2[57], oper1[61], g61[57]);
AN2 GA61_58(oper2[58], oper1[61], g61[58]);
AN2 GA61_59(oper2[59], oper1[61], g61[59]);
AN2 GA61_60(oper2[60], oper1[61], g61[60]);
AN2 GA61_61(oper2[61], oper1[61], g61[61]);
AN2 GA61_62(oper2[62], oper1[61], g61[62]);
AN2 GA61_63(oper2[63], oper1[61], g61[63]);
AN2 GA60_8(oper2[8], oper1[60], g60[8]);
AN2 GA60_9(oper2[9], oper1[60], g60[9]);
AN2 GA60_10(oper2[10], oper1[60], g60[10]);
AN2 GA60_11(oper2[11], oper1[60], g60[11]);
AN2 GA60_12(oper2[12], oper1[60], g60[12]);
AN2 GA60_13(oper2[13], oper1[60], g60[13]);
AN2 GA60_14(oper2[14], oper1[60], g60[14]);
AN2 GA60_15(oper2[15], oper1[60], g60[15]);
AN2 GA60_16(oper2[16], oper1[60], g60[16]);
AN2 GA60_17(oper2[17], oper1[60], g60[17]);
AN2 GA60_18(oper2[18], oper1[60], g60[18]);
AN2 GA60_19(oper2[19], oper1[60], g60[19]);
AN2 GA60_20(oper2[20], oper1[60], g60[20]);
AN2 GA60_21(oper2[21], oper1[60], g60[21]);
AN2 GA60_22(oper2[22], oper1[60], g60[22]);
AN2 GA60_23(oper2[23], oper1[60], g60[23]);
AN2 GA60_24(oper2[24], oper1[60], g60[24]);
AN2 GA60_25(oper2[25], oper1[60], g60[25]);
AN2 GA60_26(oper2[26], oper1[60], g60[26]);
AN2 GA60_27(oper2[27], oper1[60], g60[27]);
AN2 GA60_28(oper2[28], oper1[60], g60[28]);
AN2 GA60_29(oper2[29], oper1[60], g60[29]);
AN2 GA60_30(oper2[30], oper1[60], g60[30]);
AN2 GA60_31(oper2[31], oper1[60], g60[31]);
AN2 GA60_32(oper2[32], oper1[60], g60[32]);
AN2 GA60_33(oper2[33], oper1[60], g60[33]);
AN2 GA60_34(oper2[34], oper1[60], g60[34]);
AN2 GA60_35(oper2[35], oper1[60], g60[35]);
AN2 GA60_36(oper2[36], oper1[60], g60[36]);
AN2 GA60_37(oper2[37], oper1[60], g60[37]);
AN2 GA60_38(oper2[38], oper1[60], g60[38]);
AN2 GA60_39(oper2[39], oper1[60], g60[39]);
AN2 GA60_40(oper2[40], oper1[60], g60[40]);
AN2 GA60_41(oper2[41], oper1[60], g60[41]);
AN2 GA60_42(oper2[42], oper1[60], g60[42]);
AN2 GA60_43(oper2[43], oper1[60], g60[43]);
AN2 GA60_44(oper2[44], oper1[60], g60[44]);
AN2 GA60_45(oper2[45], oper1[60], g60[45]);
AN2 GA60_46(oper2[46], oper1[60], g60[46]);
AN2 GA60_47(oper2[47], oper1[60], g60[47]);
AN2 GA60_48(oper2[48], oper1[60], g60[48]);
AN2 GA60_49(oper2[49], oper1[60], g60[49]);
AN2 GA60_50(oper2[50], oper1[60], g60[50]);
AN2 GA60_51(oper2[51], oper1[60], g60[51]);
AN2 GA60_52(oper2[52], oper1[60], g60[52]);
AN2 GA60_53(oper2[53], oper1[60], g60[53]);
AN2 GA60_54(oper2[54], oper1[60], g60[54]);
AN2 GA60_55(oper2[55], oper1[60], g60[55]);
AN2 GA60_56(oper2[56], oper1[60], g60[56]);
AN2 GA60_57(oper2[57], oper1[60], g60[57]);
AN2 GA60_58(oper2[58], oper1[60], g60[58]);
AN2 GA60_59(oper2[59], oper1[60], g60[59]);
AN2 GA60_60(oper2[60], oper1[60], g60[60]);
AN2 GA60_61(oper2[61], oper1[60], g60[61]);
AN2 GA60_62(oper2[62], oper1[60], g60[62]);
AN2 GA60_63(oper2[63], oper1[60], g60[63]);
AN2 GA59_8(oper2[8], oper1[59], g59[8]);
AN2 GA59_9(oper2[9], oper1[59], g59[9]);
AN2 GA59_10(oper2[10], oper1[59], g59[10]);
AN2 GA59_11(oper2[11], oper1[59], g59[11]);
AN2 GA59_12(oper2[12], oper1[59], g59[12]);
AN2 GA59_13(oper2[13], oper1[59], g59[13]);
AN2 GA59_14(oper2[14], oper1[59], g59[14]);
AN2 GA59_15(oper2[15], oper1[59], g59[15]);
AN2 GA59_16(oper2[16], oper1[59], g59[16]);
AN2 GA59_17(oper2[17], oper1[59], g59[17]);
AN2 GA59_18(oper2[18], oper1[59], g59[18]);
AN2 GA59_19(oper2[19], oper1[59], g59[19]);
AN2 GA59_20(oper2[20], oper1[59], g59[20]);
AN2 GA59_21(oper2[21], oper1[59], g59[21]);
AN2 GA59_22(oper2[22], oper1[59], g59[22]);
AN2 GA59_23(oper2[23], oper1[59], g59[23]);
AN2 GA59_24(oper2[24], oper1[59], g59[24]);
AN2 GA59_25(oper2[25], oper1[59], g59[25]);
AN2 GA59_26(oper2[26], oper1[59], g59[26]);
AN2 GA59_27(oper2[27], oper1[59], g59[27]);
AN2 GA59_28(oper2[28], oper1[59], g59[28]);
AN2 GA59_29(oper2[29], oper1[59], g59[29]);
AN2 GA59_30(oper2[30], oper1[59], g59[30]);
AN2 GA59_31(oper2[31], oper1[59], g59[31]);
AN2 GA59_32(oper2[32], oper1[59], g59[32]);
AN2 GA59_33(oper2[33], oper1[59], g59[33]);
AN2 GA59_34(oper2[34], oper1[59], g59[34]);
AN2 GA59_35(oper2[35], oper1[59], g59[35]);
AN2 GA59_36(oper2[36], oper1[59], g59[36]);
AN2 GA59_37(oper2[37], oper1[59], g59[37]);
AN2 GA59_38(oper2[38], oper1[59], g59[38]);
AN2 GA59_39(oper2[39], oper1[59], g59[39]);
AN2 GA59_40(oper2[40], oper1[59], g59[40]);
AN2 GA59_41(oper2[41], oper1[59], g59[41]);
AN2 GA59_42(oper2[42], oper1[59], g59[42]);
AN2 GA59_43(oper2[43], oper1[59], g59[43]);
AN2 GA59_44(oper2[44], oper1[59], g59[44]);
AN2 GA59_45(oper2[45], oper1[59], g59[45]);
AN2 GA59_46(oper2[46], oper1[59], g59[46]);
AN2 GA59_47(oper2[47], oper1[59], g59[47]);
AN2 GA59_48(oper2[48], oper1[59], g59[48]);
AN2 GA59_49(oper2[49], oper1[59], g59[49]);
AN2 GA59_50(oper2[50], oper1[59], g59[50]);
AN2 GA59_51(oper2[51], oper1[59], g59[51]);
AN2 GA59_52(oper2[52], oper1[59], g59[52]);
AN2 GA59_53(oper2[53], oper1[59], g59[53]);
AN2 GA59_54(oper2[54], oper1[59], g59[54]);
AN2 GA59_55(oper2[55], oper1[59], g59[55]);
AN2 GA59_56(oper2[56], oper1[59], g59[56]);
AN2 GA59_57(oper2[57], oper1[59], g59[57]);
AN2 GA59_58(oper2[58], oper1[59], g59[58]);
AN2 GA59_59(oper2[59], oper1[59], g59[59]);
AN2 GA59_60(oper2[60], oper1[59], g59[60]);
AN2 GA59_61(oper2[61], oper1[59], g59[61]);
AN2 GA59_62(oper2[62], oper1[59], g59[62]);
AN2 GA59_63(oper2[63], oper1[59], g59[63]);
AN2 GA58_8(oper2[8], oper1[58], g58[8]);
AN2 GA58_9(oper2[9], oper1[58], g58[9]);
AN2 GA58_10(oper2[10], oper1[58], g58[10]);
AN2 GA58_11(oper2[11], oper1[58], g58[11]);
AN2 GA58_12(oper2[12], oper1[58], g58[12]);
AN2 GA58_13(oper2[13], oper1[58], g58[13]);
AN2 GA58_14(oper2[14], oper1[58], g58[14]);
AN2 GA58_15(oper2[15], oper1[58], g58[15]);
AN2 GA58_16(oper2[16], oper1[58], g58[16]);
AN2 GA58_17(oper2[17], oper1[58], g58[17]);
AN2 GA58_18(oper2[18], oper1[58], g58[18]);
AN2 GA58_19(oper2[19], oper1[58], g58[19]);
AN2 GA58_20(oper2[20], oper1[58], g58[20]);
AN2 GA58_21(oper2[21], oper1[58], g58[21]);
AN2 GA58_22(oper2[22], oper1[58], g58[22]);
AN2 GA58_23(oper2[23], oper1[58], g58[23]);
AN2 GA58_24(oper2[24], oper1[58], g58[24]);
AN2 GA58_25(oper2[25], oper1[58], g58[25]);
AN2 GA58_26(oper2[26], oper1[58], g58[26]);
AN2 GA58_27(oper2[27], oper1[58], g58[27]);
AN2 GA58_28(oper2[28], oper1[58], g58[28]);
AN2 GA58_29(oper2[29], oper1[58], g58[29]);
AN2 GA58_30(oper2[30], oper1[58], g58[30]);
AN2 GA58_31(oper2[31], oper1[58], g58[31]);
AN2 GA58_32(oper2[32], oper1[58], g58[32]);
AN2 GA58_33(oper2[33], oper1[58], g58[33]);
AN2 GA58_34(oper2[34], oper1[58], g58[34]);
AN2 GA58_35(oper2[35], oper1[58], g58[35]);
AN2 GA58_36(oper2[36], oper1[58], g58[36]);
AN2 GA58_37(oper2[37], oper1[58], g58[37]);
AN2 GA58_38(oper2[38], oper1[58], g58[38]);
AN2 GA58_39(oper2[39], oper1[58], g58[39]);
AN2 GA58_40(oper2[40], oper1[58], g58[40]);
AN2 GA58_41(oper2[41], oper1[58], g58[41]);
AN2 GA58_42(oper2[42], oper1[58], g58[42]);
AN2 GA58_43(oper2[43], oper1[58], g58[43]);
AN2 GA58_44(oper2[44], oper1[58], g58[44]);
AN2 GA58_45(oper2[45], oper1[58], g58[45]);
AN2 GA58_46(oper2[46], oper1[58], g58[46]);
AN2 GA58_47(oper2[47], oper1[58], g58[47]);
AN2 GA58_48(oper2[48], oper1[58], g58[48]);
AN2 GA58_49(oper2[49], oper1[58], g58[49]);
AN2 GA58_50(oper2[50], oper1[58], g58[50]);
AN2 GA58_51(oper2[51], oper1[58], g58[51]);
AN2 GA58_52(oper2[52], oper1[58], g58[52]);
AN2 GA58_53(oper2[53], oper1[58], g58[53]);
AN2 GA58_54(oper2[54], oper1[58], g58[54]);
AN2 GA58_55(oper2[55], oper1[58], g58[55]);
AN2 GA58_56(oper2[56], oper1[58], g58[56]);
AN2 GA58_57(oper2[57], oper1[58], g58[57]);
AN2 GA58_58(oper2[58], oper1[58], g58[58]);
AN2 GA58_59(oper2[59], oper1[58], g58[59]);
AN2 GA58_60(oper2[60], oper1[58], g58[60]);
AN2 GA58_61(oper2[61], oper1[58], g58[61]);
AN2 GA58_62(oper2[62], oper1[58], g58[62]);
AN2 GA58_63(oper2[63], oper1[58], g58[63]);
AN2 GA57_8(oper2[8], oper1[57], g57[8]);
AN2 GA57_9(oper2[9], oper1[57], g57[9]);
AN2 GA57_10(oper2[10], oper1[57], g57[10]);
AN2 GA57_11(oper2[11], oper1[57], g57[11]);
AN2 GA57_12(oper2[12], oper1[57], g57[12]);
AN2 GA57_13(oper2[13], oper1[57], g57[13]);
AN2 GA57_14(oper2[14], oper1[57], g57[14]);
AN2 GA57_15(oper2[15], oper1[57], g57[15]);
AN2 GA57_16(oper2[16], oper1[57], g57[16]);
AN2 GA57_17(oper2[17], oper1[57], g57[17]);
AN2 GA57_18(oper2[18], oper1[57], g57[18]);
AN2 GA57_19(oper2[19], oper1[57], g57[19]);
AN2 GA57_20(oper2[20], oper1[57], g57[20]);
AN2 GA57_21(oper2[21], oper1[57], g57[21]);
AN2 GA57_22(oper2[22], oper1[57], g57[22]);
AN2 GA57_23(oper2[23], oper1[57], g57[23]);
AN2 GA57_24(oper2[24], oper1[57], g57[24]);
AN2 GA57_25(oper2[25], oper1[57], g57[25]);
AN2 GA57_26(oper2[26], oper1[57], g57[26]);
AN2 GA57_27(oper2[27], oper1[57], g57[27]);
AN2 GA57_28(oper2[28], oper1[57], g57[28]);
AN2 GA57_29(oper2[29], oper1[57], g57[29]);
AN2 GA57_30(oper2[30], oper1[57], g57[30]);
AN2 GA57_31(oper2[31], oper1[57], g57[31]);
AN2 GA57_32(oper2[32], oper1[57], g57[32]);
AN2 GA57_33(oper2[33], oper1[57], g57[33]);
AN2 GA57_34(oper2[34], oper1[57], g57[34]);
AN2 GA57_35(oper2[35], oper1[57], g57[35]);
AN2 GA57_36(oper2[36], oper1[57], g57[36]);
AN2 GA57_37(oper2[37], oper1[57], g57[37]);
AN2 GA57_38(oper2[38], oper1[57], g57[38]);
AN2 GA57_39(oper2[39], oper1[57], g57[39]);
AN2 GA57_40(oper2[40], oper1[57], g57[40]);
AN2 GA57_41(oper2[41], oper1[57], g57[41]);
AN2 GA57_42(oper2[42], oper1[57], g57[42]);
AN2 GA57_43(oper2[43], oper1[57], g57[43]);
AN2 GA57_44(oper2[44], oper1[57], g57[44]);
AN2 GA57_45(oper2[45], oper1[57], g57[45]);
AN2 GA57_46(oper2[46], oper1[57], g57[46]);
AN2 GA57_47(oper2[47], oper1[57], g57[47]);
AN2 GA57_48(oper2[48], oper1[57], g57[48]);
AN2 GA57_49(oper2[49], oper1[57], g57[49]);
AN2 GA57_50(oper2[50], oper1[57], g57[50]);
AN2 GA57_51(oper2[51], oper1[57], g57[51]);
AN2 GA57_52(oper2[52], oper1[57], g57[52]);
AN2 GA57_53(oper2[53], oper1[57], g57[53]);
AN2 GA57_54(oper2[54], oper1[57], g57[54]);
AN2 GA57_55(oper2[55], oper1[57], g57[55]);
AN2 GA57_56(oper2[56], oper1[57], g57[56]);
AN2 GA57_57(oper2[57], oper1[57], g57[57]);
AN2 GA57_58(oper2[58], oper1[57], g57[58]);
AN2 GA57_59(oper2[59], oper1[57], g57[59]);
AN2 GA57_60(oper2[60], oper1[57], g57[60]);
AN2 GA57_61(oper2[61], oper1[57], g57[61]);
AN2 GA57_62(oper2[62], oper1[57], g57[62]);
AN2 GA57_63(oper2[63], oper1[57], g57[63]);
AN2 GA56_8(oper2[8], oper1[56], g56[8]);
AN2 GA56_9(oper2[9], oper1[56], g56[9]);
AN2 GA56_10(oper2[10], oper1[56], g56[10]);
AN2 GA56_11(oper2[11], oper1[56], g56[11]);
AN2 GA56_12(oper2[12], oper1[56], g56[12]);
AN2 GA56_13(oper2[13], oper1[56], g56[13]);
AN2 GA56_14(oper2[14], oper1[56], g56[14]);
AN2 GA56_15(oper2[15], oper1[56], g56[15]);
AN2 GA56_16(oper2[16], oper1[56], g56[16]);
AN2 GA56_17(oper2[17], oper1[56], g56[17]);
AN2 GA56_18(oper2[18], oper1[56], g56[18]);
AN2 GA56_19(oper2[19], oper1[56], g56[19]);
AN2 GA56_20(oper2[20], oper1[56], g56[20]);
AN2 GA56_21(oper2[21], oper1[56], g56[21]);
AN2 GA56_22(oper2[22], oper1[56], g56[22]);
AN2 GA56_23(oper2[23], oper1[56], g56[23]);
AN2 GA56_24(oper2[24], oper1[56], g56[24]);
AN2 GA56_25(oper2[25], oper1[56], g56[25]);
AN2 GA56_26(oper2[26], oper1[56], g56[26]);
AN2 GA56_27(oper2[27], oper1[56], g56[27]);
AN2 GA56_28(oper2[28], oper1[56], g56[28]);
AN2 GA56_29(oper2[29], oper1[56], g56[29]);
AN2 GA56_30(oper2[30], oper1[56], g56[30]);
AN2 GA56_31(oper2[31], oper1[56], g56[31]);
AN2 GA56_32(oper2[32], oper1[56], g56[32]);
AN2 GA56_33(oper2[33], oper1[56], g56[33]);
AN2 GA56_34(oper2[34], oper1[56], g56[34]);
AN2 GA56_35(oper2[35], oper1[56], g56[35]);
AN2 GA56_36(oper2[36], oper1[56], g56[36]);
AN2 GA56_37(oper2[37], oper1[56], g56[37]);
AN2 GA56_38(oper2[38], oper1[56], g56[38]);
AN2 GA56_39(oper2[39], oper1[56], g56[39]);
AN2 GA56_40(oper2[40], oper1[56], g56[40]);
AN2 GA56_41(oper2[41], oper1[56], g56[41]);
AN2 GA56_42(oper2[42], oper1[56], g56[42]);
AN2 GA56_43(oper2[43], oper1[56], g56[43]);
AN2 GA56_44(oper2[44], oper1[56], g56[44]);
AN2 GA56_45(oper2[45], oper1[56], g56[45]);
AN2 GA56_46(oper2[46], oper1[56], g56[46]);
AN2 GA56_47(oper2[47], oper1[56], g56[47]);
AN2 GA56_48(oper2[48], oper1[56], g56[48]);
AN2 GA56_49(oper2[49], oper1[56], g56[49]);
AN2 GA56_50(oper2[50], oper1[56], g56[50]);
AN2 GA56_51(oper2[51], oper1[56], g56[51]);
AN2 GA56_52(oper2[52], oper1[56], g56[52]);
AN2 GA56_53(oper2[53], oper1[56], g56[53]);
AN2 GA56_54(oper2[54], oper1[56], g56[54]);
AN2 GA56_55(oper2[55], oper1[56], g56[55]);
AN2 GA56_56(oper2[56], oper1[56], g56[56]);
AN2 GA56_57(oper2[57], oper1[56], g56[57]);
AN2 GA56_58(oper2[58], oper1[56], g56[58]);
AN2 GA56_59(oper2[59], oper1[56], g56[59]);
AN2 GA56_60(oper2[60], oper1[56], g56[60]);
AN2 GA56_61(oper2[61], oper1[56], g56[61]);
AN2 GA56_62(oper2[62], oper1[56], g56[62]);
AN2 GA56_63(oper2[63], oper1[56], g56[63]);
AN2 GA55_8(oper2[8], oper1[55], g55[8]);
AN2 GA55_9(oper2[9], oper1[55], g55[9]);
AN2 GA55_10(oper2[10], oper1[55], g55[10]);
AN2 GA55_11(oper2[11], oper1[55], g55[11]);
AN2 GA55_12(oper2[12], oper1[55], g55[12]);
AN2 GA55_13(oper2[13], oper1[55], g55[13]);
AN2 GA55_14(oper2[14], oper1[55], g55[14]);
AN2 GA55_15(oper2[15], oper1[55], g55[15]);
AN2 GA55_16(oper2[16], oper1[55], g55[16]);
AN2 GA55_17(oper2[17], oper1[55], g55[17]);
AN2 GA55_18(oper2[18], oper1[55], g55[18]);
AN2 GA55_19(oper2[19], oper1[55], g55[19]);
AN2 GA55_20(oper2[20], oper1[55], g55[20]);
AN2 GA55_21(oper2[21], oper1[55], g55[21]);
AN2 GA55_22(oper2[22], oper1[55], g55[22]);
AN2 GA55_23(oper2[23], oper1[55], g55[23]);
AN2 GA55_24(oper2[24], oper1[55], g55[24]);
AN2 GA55_25(oper2[25], oper1[55], g55[25]);
AN2 GA55_26(oper2[26], oper1[55], g55[26]);
AN2 GA55_27(oper2[27], oper1[55], g55[27]);
AN2 GA55_28(oper2[28], oper1[55], g55[28]);
AN2 GA55_29(oper2[29], oper1[55], g55[29]);
AN2 GA55_30(oper2[30], oper1[55], g55[30]);
AN2 GA55_31(oper2[31], oper1[55], g55[31]);
AN2 GA55_32(oper2[32], oper1[55], g55[32]);
AN2 GA55_33(oper2[33], oper1[55], g55[33]);
AN2 GA55_34(oper2[34], oper1[55], g55[34]);
AN2 GA55_35(oper2[35], oper1[55], g55[35]);
AN2 GA55_36(oper2[36], oper1[55], g55[36]);
AN2 GA55_37(oper2[37], oper1[55], g55[37]);
AN2 GA55_38(oper2[38], oper1[55], g55[38]);
AN2 GA55_39(oper2[39], oper1[55], g55[39]);
AN2 GA55_40(oper2[40], oper1[55], g55[40]);
AN2 GA55_41(oper2[41], oper1[55], g55[41]);
AN2 GA55_42(oper2[42], oper1[55], g55[42]);
AN2 GA55_43(oper2[43], oper1[55], g55[43]);
AN2 GA55_44(oper2[44], oper1[55], g55[44]);
AN2 GA55_45(oper2[45], oper1[55], g55[45]);
AN2 GA55_46(oper2[46], oper1[55], g55[46]);
AN2 GA55_47(oper2[47], oper1[55], g55[47]);
AN2 GA55_48(oper2[48], oper1[55], g55[48]);
AN2 GA55_49(oper2[49], oper1[55], g55[49]);
AN2 GA55_50(oper2[50], oper1[55], g55[50]);
AN2 GA55_51(oper2[51], oper1[55], g55[51]);
AN2 GA55_52(oper2[52], oper1[55], g55[52]);
AN2 GA55_53(oper2[53], oper1[55], g55[53]);
AN2 GA55_54(oper2[54], oper1[55], g55[54]);
AN2 GA55_55(oper2[55], oper1[55], g55[55]);
AN2 GA55_56(oper2[56], oper1[55], g55[56]);
AN2 GA55_57(oper2[57], oper1[55], g55[57]);
AN2 GA55_58(oper2[58], oper1[55], g55[58]);
AN2 GA55_59(oper2[59], oper1[55], g55[59]);
AN2 GA55_60(oper2[60], oper1[55], g55[60]);
AN2 GA55_61(oper2[61], oper1[55], g55[61]);
AN2 GA55_62(oper2[62], oper1[55], g55[62]);
AN2 GA55_63(oper2[63], oper1[55], g55[63]);
AN2 GA54_8(oper2[8], oper1[54], g54[8]);
AN2 GA54_9(oper2[9], oper1[54], g54[9]);
AN2 GA54_10(oper2[10], oper1[54], g54[10]);
AN2 GA54_11(oper2[11], oper1[54], g54[11]);
AN2 GA54_12(oper2[12], oper1[54], g54[12]);
AN2 GA54_13(oper2[13], oper1[54], g54[13]);
AN2 GA54_14(oper2[14], oper1[54], g54[14]);
AN2 GA54_15(oper2[15], oper1[54], g54[15]);
AN2 GA54_16(oper2[16], oper1[54], g54[16]);
AN2 GA54_17(oper2[17], oper1[54], g54[17]);
AN2 GA54_18(oper2[18], oper1[54], g54[18]);
AN2 GA54_19(oper2[19], oper1[54], g54[19]);
AN2 GA54_20(oper2[20], oper1[54], g54[20]);
AN2 GA54_21(oper2[21], oper1[54], g54[21]);
AN2 GA54_22(oper2[22], oper1[54], g54[22]);
AN2 GA54_23(oper2[23], oper1[54], g54[23]);
AN2 GA54_24(oper2[24], oper1[54], g54[24]);
AN2 GA54_25(oper2[25], oper1[54], g54[25]);
AN2 GA54_26(oper2[26], oper1[54], g54[26]);
AN2 GA54_27(oper2[27], oper1[54], g54[27]);
AN2 GA54_28(oper2[28], oper1[54], g54[28]);
AN2 GA54_29(oper2[29], oper1[54], g54[29]);
AN2 GA54_30(oper2[30], oper1[54], g54[30]);
AN2 GA54_31(oper2[31], oper1[54], g54[31]);
AN2 GA54_32(oper2[32], oper1[54], g54[32]);
AN2 GA54_33(oper2[33], oper1[54], g54[33]);
AN2 GA54_34(oper2[34], oper1[54], g54[34]);
AN2 GA54_35(oper2[35], oper1[54], g54[35]);
AN2 GA54_36(oper2[36], oper1[54], g54[36]);
AN2 GA54_37(oper2[37], oper1[54], g54[37]);
AN2 GA54_38(oper2[38], oper1[54], g54[38]);
AN2 GA54_39(oper2[39], oper1[54], g54[39]);
AN2 GA54_40(oper2[40], oper1[54], g54[40]);
AN2 GA54_41(oper2[41], oper1[54], g54[41]);
AN2 GA54_42(oper2[42], oper1[54], g54[42]);
AN2 GA54_43(oper2[43], oper1[54], g54[43]);
AN2 GA54_44(oper2[44], oper1[54], g54[44]);
AN2 GA54_45(oper2[45], oper1[54], g54[45]);
AN2 GA54_46(oper2[46], oper1[54], g54[46]);
AN2 GA54_47(oper2[47], oper1[54], g54[47]);
AN2 GA54_48(oper2[48], oper1[54], g54[48]);
AN2 GA54_49(oper2[49], oper1[54], g54[49]);
AN2 GA54_50(oper2[50], oper1[54], g54[50]);
AN2 GA54_51(oper2[51], oper1[54], g54[51]);
AN2 GA54_52(oper2[52], oper1[54], g54[52]);
AN2 GA54_53(oper2[53], oper1[54], g54[53]);
AN2 GA54_54(oper2[54], oper1[54], g54[54]);
AN2 GA54_55(oper2[55], oper1[54], g54[55]);
AN2 GA54_56(oper2[56], oper1[54], g54[56]);
AN2 GA54_57(oper2[57], oper1[54], g54[57]);
AN2 GA54_58(oper2[58], oper1[54], g54[58]);
AN2 GA54_59(oper2[59], oper1[54], g54[59]);
AN2 GA54_60(oper2[60], oper1[54], g54[60]);
AN2 GA54_61(oper2[61], oper1[54], g54[61]);
AN2 GA54_62(oper2[62], oper1[54], g54[62]);
AN2 GA54_63(oper2[63], oper1[54], g54[63]);
AN2 GA53_8(oper2[8], oper1[53], g53[8]);
AN2 GA53_9(oper2[9], oper1[53], g53[9]);
AN2 GA53_10(oper2[10], oper1[53], g53[10]);
AN2 GA53_11(oper2[11], oper1[53], g53[11]);
AN2 GA53_12(oper2[12], oper1[53], g53[12]);
AN2 GA53_13(oper2[13], oper1[53], g53[13]);
AN2 GA53_14(oper2[14], oper1[53], g53[14]);
AN2 GA53_15(oper2[15], oper1[53], g53[15]);
AN2 GA53_16(oper2[16], oper1[53], g53[16]);
AN2 GA53_17(oper2[17], oper1[53], g53[17]);
AN2 GA53_18(oper2[18], oper1[53], g53[18]);
AN2 GA53_19(oper2[19], oper1[53], g53[19]);
AN2 GA53_20(oper2[20], oper1[53], g53[20]);
AN2 GA53_21(oper2[21], oper1[53], g53[21]);
AN2 GA53_22(oper2[22], oper1[53], g53[22]);
AN2 GA53_23(oper2[23], oper1[53], g53[23]);
AN2 GA53_24(oper2[24], oper1[53], g53[24]);
AN2 GA53_25(oper2[25], oper1[53], g53[25]);
AN2 GA53_26(oper2[26], oper1[53], g53[26]);
AN2 GA53_27(oper2[27], oper1[53], g53[27]);
AN2 GA53_28(oper2[28], oper1[53], g53[28]);
AN2 GA53_29(oper2[29], oper1[53], g53[29]);
AN2 GA53_30(oper2[30], oper1[53], g53[30]);
AN2 GA53_31(oper2[31], oper1[53], g53[31]);
AN2 GA53_32(oper2[32], oper1[53], g53[32]);
AN2 GA53_33(oper2[33], oper1[53], g53[33]);
AN2 GA53_34(oper2[34], oper1[53], g53[34]);
AN2 GA53_35(oper2[35], oper1[53], g53[35]);
AN2 GA53_36(oper2[36], oper1[53], g53[36]);
AN2 GA53_37(oper2[37], oper1[53], g53[37]);
AN2 GA53_38(oper2[38], oper1[53], g53[38]);
AN2 GA53_39(oper2[39], oper1[53], g53[39]);
AN2 GA53_40(oper2[40], oper1[53], g53[40]);
AN2 GA53_41(oper2[41], oper1[53], g53[41]);
AN2 GA53_42(oper2[42], oper1[53], g53[42]);
AN2 GA53_43(oper2[43], oper1[53], g53[43]);
AN2 GA53_44(oper2[44], oper1[53], g53[44]);
AN2 GA53_45(oper2[45], oper1[53], g53[45]);
AN2 GA53_46(oper2[46], oper1[53], g53[46]);
AN2 GA53_47(oper2[47], oper1[53], g53[47]);
AN2 GA53_48(oper2[48], oper1[53], g53[48]);
AN2 GA53_49(oper2[49], oper1[53], g53[49]);
AN2 GA53_50(oper2[50], oper1[53], g53[50]);
AN2 GA53_51(oper2[51], oper1[53], g53[51]);
AN2 GA53_52(oper2[52], oper1[53], g53[52]);
AN2 GA53_53(oper2[53], oper1[53], g53[53]);
AN2 GA53_54(oper2[54], oper1[53], g53[54]);
AN2 GA53_55(oper2[55], oper1[53], g53[55]);
AN2 GA53_56(oper2[56], oper1[53], g53[56]);
AN2 GA53_57(oper2[57], oper1[53], g53[57]);
AN2 GA53_58(oper2[58], oper1[53], g53[58]);
AN2 GA53_59(oper2[59], oper1[53], g53[59]);
AN2 GA53_60(oper2[60], oper1[53], g53[60]);
AN2 GA53_61(oper2[61], oper1[53], g53[61]);
AN2 GA53_62(oper2[62], oper1[53], g53[62]);
AN2 GA53_63(oper2[63], oper1[53], g53[63]);
AN2 GA52_8(oper2[8], oper1[52], g52[8]);
AN2 GA52_9(oper2[9], oper1[52], g52[9]);
AN2 GA52_10(oper2[10], oper1[52], g52[10]);
AN2 GA52_11(oper2[11], oper1[52], g52[11]);
AN2 GA52_12(oper2[12], oper1[52], g52[12]);
AN2 GA52_13(oper2[13], oper1[52], g52[13]);
AN2 GA52_14(oper2[14], oper1[52], g52[14]);
AN2 GA52_15(oper2[15], oper1[52], g52[15]);
AN2 GA52_16(oper2[16], oper1[52], g52[16]);
AN2 GA52_17(oper2[17], oper1[52], g52[17]);
AN2 GA52_18(oper2[18], oper1[52], g52[18]);
AN2 GA52_19(oper2[19], oper1[52], g52[19]);
AN2 GA52_20(oper2[20], oper1[52], g52[20]);
AN2 GA52_21(oper2[21], oper1[52], g52[21]);
AN2 GA52_22(oper2[22], oper1[52], g52[22]);
AN2 GA52_23(oper2[23], oper1[52], g52[23]);
AN2 GA52_24(oper2[24], oper1[52], g52[24]);
AN2 GA52_25(oper2[25], oper1[52], g52[25]);
AN2 GA52_26(oper2[26], oper1[52], g52[26]);
AN2 GA52_27(oper2[27], oper1[52], g52[27]);
AN2 GA52_28(oper2[28], oper1[52], g52[28]);
AN2 GA52_29(oper2[29], oper1[52], g52[29]);
AN2 GA52_30(oper2[30], oper1[52], g52[30]);
AN2 GA52_31(oper2[31], oper1[52], g52[31]);
AN2 GA52_32(oper2[32], oper1[52], g52[32]);
AN2 GA52_33(oper2[33], oper1[52], g52[33]);
AN2 GA52_34(oper2[34], oper1[52], g52[34]);
AN2 GA52_35(oper2[35], oper1[52], g52[35]);
AN2 GA52_36(oper2[36], oper1[52], g52[36]);
AN2 GA52_37(oper2[37], oper1[52], g52[37]);
AN2 GA52_38(oper2[38], oper1[52], g52[38]);
AN2 GA52_39(oper2[39], oper1[52], g52[39]);
AN2 GA52_40(oper2[40], oper1[52], g52[40]);
AN2 GA52_41(oper2[41], oper1[52], g52[41]);
AN2 GA52_42(oper2[42], oper1[52], g52[42]);
AN2 GA52_43(oper2[43], oper1[52], g52[43]);
AN2 GA52_44(oper2[44], oper1[52], g52[44]);
AN2 GA52_45(oper2[45], oper1[52], g52[45]);
AN2 GA52_46(oper2[46], oper1[52], g52[46]);
AN2 GA52_47(oper2[47], oper1[52], g52[47]);
AN2 GA52_48(oper2[48], oper1[52], g52[48]);
AN2 GA52_49(oper2[49], oper1[52], g52[49]);
AN2 GA52_50(oper2[50], oper1[52], g52[50]);
AN2 GA52_51(oper2[51], oper1[52], g52[51]);
AN2 GA52_52(oper2[52], oper1[52], g52[52]);
AN2 GA52_53(oper2[53], oper1[52], g52[53]);
AN2 GA52_54(oper2[54], oper1[52], g52[54]);
AN2 GA52_55(oper2[55], oper1[52], g52[55]);
AN2 GA52_56(oper2[56], oper1[52], g52[56]);
AN2 GA52_57(oper2[57], oper1[52], g52[57]);
AN2 GA52_58(oper2[58], oper1[52], g52[58]);
AN2 GA52_59(oper2[59], oper1[52], g52[59]);
AN2 GA52_60(oper2[60], oper1[52], g52[60]);
AN2 GA52_61(oper2[61], oper1[52], g52[61]);
AN2 GA52_62(oper2[62], oper1[52], g52[62]);
AN2 GA52_63(oper2[63], oper1[52], g52[63]);
AN2 GA51_8(oper2[8], oper1[51], g51[8]);
AN2 GA51_9(oper2[9], oper1[51], g51[9]);
AN2 GA51_10(oper2[10], oper1[51], g51[10]);
AN2 GA51_11(oper2[11], oper1[51], g51[11]);
AN2 GA51_12(oper2[12], oper1[51], g51[12]);
AN2 GA51_13(oper2[13], oper1[51], g51[13]);
AN2 GA51_14(oper2[14], oper1[51], g51[14]);
AN2 GA51_15(oper2[15], oper1[51], g51[15]);
AN2 GA51_16(oper2[16], oper1[51], g51[16]);
AN2 GA51_17(oper2[17], oper1[51], g51[17]);
AN2 GA51_18(oper2[18], oper1[51], g51[18]);
AN2 GA51_19(oper2[19], oper1[51], g51[19]);
AN2 GA51_20(oper2[20], oper1[51], g51[20]);
AN2 GA51_21(oper2[21], oper1[51], g51[21]);
AN2 GA51_22(oper2[22], oper1[51], g51[22]);
AN2 GA51_23(oper2[23], oper1[51], g51[23]);
AN2 GA51_24(oper2[24], oper1[51], g51[24]);
AN2 GA51_25(oper2[25], oper1[51], g51[25]);
AN2 GA51_26(oper2[26], oper1[51], g51[26]);
AN2 GA51_27(oper2[27], oper1[51], g51[27]);
AN2 GA51_28(oper2[28], oper1[51], g51[28]);
AN2 GA51_29(oper2[29], oper1[51], g51[29]);
AN2 GA51_30(oper2[30], oper1[51], g51[30]);
AN2 GA51_31(oper2[31], oper1[51], g51[31]);
AN2 GA51_32(oper2[32], oper1[51], g51[32]);
AN2 GA51_33(oper2[33], oper1[51], g51[33]);
AN2 GA51_34(oper2[34], oper1[51], g51[34]);
AN2 GA51_35(oper2[35], oper1[51], g51[35]);
AN2 GA51_36(oper2[36], oper1[51], g51[36]);
AN2 GA51_37(oper2[37], oper1[51], g51[37]);
AN2 GA51_38(oper2[38], oper1[51], g51[38]);
AN2 GA51_39(oper2[39], oper1[51], g51[39]);
AN2 GA51_40(oper2[40], oper1[51], g51[40]);
AN2 GA51_41(oper2[41], oper1[51], g51[41]);
AN2 GA51_42(oper2[42], oper1[51], g51[42]);
AN2 GA51_43(oper2[43], oper1[51], g51[43]);
AN2 GA51_44(oper2[44], oper1[51], g51[44]);
AN2 GA51_45(oper2[45], oper1[51], g51[45]);
AN2 GA51_46(oper2[46], oper1[51], g51[46]);
AN2 GA51_47(oper2[47], oper1[51], g51[47]);
AN2 GA51_48(oper2[48], oper1[51], g51[48]);
AN2 GA51_49(oper2[49], oper1[51], g51[49]);
AN2 GA51_50(oper2[50], oper1[51], g51[50]);
AN2 GA51_51(oper2[51], oper1[51], g51[51]);
AN2 GA51_52(oper2[52], oper1[51], g51[52]);
AN2 GA51_53(oper2[53], oper1[51], g51[53]);
AN2 GA51_54(oper2[54], oper1[51], g51[54]);
AN2 GA51_55(oper2[55], oper1[51], g51[55]);
AN2 GA51_56(oper2[56], oper1[51], g51[56]);
AN2 GA51_57(oper2[57], oper1[51], g51[57]);
AN2 GA51_58(oper2[58], oper1[51], g51[58]);
AN2 GA51_59(oper2[59], oper1[51], g51[59]);
AN2 GA51_60(oper2[60], oper1[51], g51[60]);
AN2 GA51_61(oper2[61], oper1[51], g51[61]);
AN2 GA51_62(oper2[62], oper1[51], g51[62]);
AN2 GA51_63(oper2[63], oper1[51], g51[63]);
AN2 GA50_8(oper2[8], oper1[50], g50[8]);
AN2 GA50_9(oper2[9], oper1[50], g50[9]);
AN2 GA50_10(oper2[10], oper1[50], g50[10]);
AN2 GA50_11(oper2[11], oper1[50], g50[11]);
AN2 GA50_12(oper2[12], oper1[50], g50[12]);
AN2 GA50_13(oper2[13], oper1[50], g50[13]);
AN2 GA50_14(oper2[14], oper1[50], g50[14]);
AN2 GA50_15(oper2[15], oper1[50], g50[15]);
AN2 GA50_16(oper2[16], oper1[50], g50[16]);
AN2 GA50_17(oper2[17], oper1[50], g50[17]);
AN2 GA50_18(oper2[18], oper1[50], g50[18]);
AN2 GA50_19(oper2[19], oper1[50], g50[19]);
AN2 GA50_20(oper2[20], oper1[50], g50[20]);
AN2 GA50_21(oper2[21], oper1[50], g50[21]);
AN2 GA50_22(oper2[22], oper1[50], g50[22]);
AN2 GA50_23(oper2[23], oper1[50], g50[23]);
AN2 GA50_24(oper2[24], oper1[50], g50[24]);
AN2 GA50_25(oper2[25], oper1[50], g50[25]);
AN2 GA50_26(oper2[26], oper1[50], g50[26]);
AN2 GA50_27(oper2[27], oper1[50], g50[27]);
AN2 GA50_28(oper2[28], oper1[50], g50[28]);
AN2 GA50_29(oper2[29], oper1[50], g50[29]);
AN2 GA50_30(oper2[30], oper1[50], g50[30]);
AN2 GA50_31(oper2[31], oper1[50], g50[31]);
AN2 GA50_32(oper2[32], oper1[50], g50[32]);
AN2 GA50_33(oper2[33], oper1[50], g50[33]);
AN2 GA50_34(oper2[34], oper1[50], g50[34]);
AN2 GA50_35(oper2[35], oper1[50], g50[35]);
AN2 GA50_36(oper2[36], oper1[50], g50[36]);
AN2 GA50_37(oper2[37], oper1[50], g50[37]);
AN2 GA50_38(oper2[38], oper1[50], g50[38]);
AN2 GA50_39(oper2[39], oper1[50], g50[39]);
AN2 GA50_40(oper2[40], oper1[50], g50[40]);
AN2 GA50_41(oper2[41], oper1[50], g50[41]);
AN2 GA50_42(oper2[42], oper1[50], g50[42]);
AN2 GA50_43(oper2[43], oper1[50], g50[43]);
AN2 GA50_44(oper2[44], oper1[50], g50[44]);
AN2 GA50_45(oper2[45], oper1[50], g50[45]);
AN2 GA50_46(oper2[46], oper1[50], g50[46]);
AN2 GA50_47(oper2[47], oper1[50], g50[47]);
AN2 GA50_48(oper2[48], oper1[50], g50[48]);
AN2 GA50_49(oper2[49], oper1[50], g50[49]);
AN2 GA50_50(oper2[50], oper1[50], g50[50]);
AN2 GA50_51(oper2[51], oper1[50], g50[51]);
AN2 GA50_52(oper2[52], oper1[50], g50[52]);
AN2 GA50_53(oper2[53], oper1[50], g50[53]);
AN2 GA50_54(oper2[54], oper1[50], g50[54]);
AN2 GA50_55(oper2[55], oper1[50], g50[55]);
AN2 GA50_56(oper2[56], oper1[50], g50[56]);
AN2 GA50_57(oper2[57], oper1[50], g50[57]);
AN2 GA50_58(oper2[58], oper1[50], g50[58]);
AN2 GA50_59(oper2[59], oper1[50], g50[59]);
AN2 GA50_60(oper2[60], oper1[50], g50[60]);
AN2 GA50_61(oper2[61], oper1[50], g50[61]);
AN2 GA50_62(oper2[62], oper1[50], g50[62]);
AN2 GA50_63(oper2[63], oper1[50], g50[63]);
AN2 GA49_8(oper2[8], oper1[49], g49[8]);
AN2 GA49_9(oper2[9], oper1[49], g49[9]);
AN2 GA49_10(oper2[10], oper1[49], g49[10]);
AN2 GA49_11(oper2[11], oper1[49], g49[11]);
AN2 GA49_12(oper2[12], oper1[49], g49[12]);
AN2 GA49_13(oper2[13], oper1[49], g49[13]);
AN2 GA49_14(oper2[14], oper1[49], g49[14]);
AN2 GA49_15(oper2[15], oper1[49], g49[15]);
AN2 GA49_16(oper2[16], oper1[49], g49[16]);
AN2 GA49_17(oper2[17], oper1[49], g49[17]);
AN2 GA49_18(oper2[18], oper1[49], g49[18]);
AN2 GA49_19(oper2[19], oper1[49], g49[19]);
AN2 GA49_20(oper2[20], oper1[49], g49[20]);
AN2 GA49_21(oper2[21], oper1[49], g49[21]);
AN2 GA49_22(oper2[22], oper1[49], g49[22]);
AN2 GA49_23(oper2[23], oper1[49], g49[23]);
AN2 GA49_24(oper2[24], oper1[49], g49[24]);
AN2 GA49_25(oper2[25], oper1[49], g49[25]);
AN2 GA49_26(oper2[26], oper1[49], g49[26]);
AN2 GA49_27(oper2[27], oper1[49], g49[27]);
AN2 GA49_28(oper2[28], oper1[49], g49[28]);
AN2 GA49_29(oper2[29], oper1[49], g49[29]);
AN2 GA49_30(oper2[30], oper1[49], g49[30]);
AN2 GA49_31(oper2[31], oper1[49], g49[31]);
AN2 GA49_32(oper2[32], oper1[49], g49[32]);
AN2 GA49_33(oper2[33], oper1[49], g49[33]);
AN2 GA49_34(oper2[34], oper1[49], g49[34]);
AN2 GA49_35(oper2[35], oper1[49], g49[35]);
AN2 GA49_36(oper2[36], oper1[49], g49[36]);
AN2 GA49_37(oper2[37], oper1[49], g49[37]);
AN2 GA49_38(oper2[38], oper1[49], g49[38]);
AN2 GA49_39(oper2[39], oper1[49], g49[39]);
AN2 GA49_40(oper2[40], oper1[49], g49[40]);
AN2 GA49_41(oper2[41], oper1[49], g49[41]);
AN2 GA49_42(oper2[42], oper1[49], g49[42]);
AN2 GA49_43(oper2[43], oper1[49], g49[43]);
AN2 GA49_44(oper2[44], oper1[49], g49[44]);
AN2 GA49_45(oper2[45], oper1[49], g49[45]);
AN2 GA49_46(oper2[46], oper1[49], g49[46]);
AN2 GA49_47(oper2[47], oper1[49], g49[47]);
AN2 GA49_48(oper2[48], oper1[49], g49[48]);
AN2 GA49_49(oper2[49], oper1[49], g49[49]);
AN2 GA49_50(oper2[50], oper1[49], g49[50]);
AN2 GA49_51(oper2[51], oper1[49], g49[51]);
AN2 GA49_52(oper2[52], oper1[49], g49[52]);
AN2 GA49_53(oper2[53], oper1[49], g49[53]);
AN2 GA49_54(oper2[54], oper1[49], g49[54]);
AN2 GA49_55(oper2[55], oper1[49], g49[55]);
AN2 GA49_56(oper2[56], oper1[49], g49[56]);
AN2 GA49_57(oper2[57], oper1[49], g49[57]);
AN2 GA49_58(oper2[58], oper1[49], g49[58]);
AN2 GA49_59(oper2[59], oper1[49], g49[59]);
AN2 GA49_60(oper2[60], oper1[49], g49[60]);
AN2 GA49_61(oper2[61], oper1[49], g49[61]);
AN2 GA49_62(oper2[62], oper1[49], g49[62]);
AN2 GA49_63(oper2[63], oper1[49], g49[63]);
AN2 GA48_8(oper2[8], oper1[48], g48[8]);
AN2 GA48_9(oper2[9], oper1[48], g48[9]);
AN2 GA48_10(oper2[10], oper1[48], g48[10]);
AN2 GA48_11(oper2[11], oper1[48], g48[11]);
AN2 GA48_12(oper2[12], oper1[48], g48[12]);
AN2 GA48_13(oper2[13], oper1[48], g48[13]);
AN2 GA48_14(oper2[14], oper1[48], g48[14]);
AN2 GA48_15(oper2[15], oper1[48], g48[15]);
AN2 GA48_16(oper2[16], oper1[48], g48[16]);
AN2 GA48_17(oper2[17], oper1[48], g48[17]);
AN2 GA48_18(oper2[18], oper1[48], g48[18]);
AN2 GA48_19(oper2[19], oper1[48], g48[19]);
AN2 GA48_20(oper2[20], oper1[48], g48[20]);
AN2 GA48_21(oper2[21], oper1[48], g48[21]);
AN2 GA48_22(oper2[22], oper1[48], g48[22]);
AN2 GA48_23(oper2[23], oper1[48], g48[23]);
AN2 GA48_24(oper2[24], oper1[48], g48[24]);
AN2 GA48_25(oper2[25], oper1[48], g48[25]);
AN2 GA48_26(oper2[26], oper1[48], g48[26]);
AN2 GA48_27(oper2[27], oper1[48], g48[27]);
AN2 GA48_28(oper2[28], oper1[48], g48[28]);
AN2 GA48_29(oper2[29], oper1[48], g48[29]);
AN2 GA48_30(oper2[30], oper1[48], g48[30]);
AN2 GA48_31(oper2[31], oper1[48], g48[31]);
AN2 GA48_32(oper2[32], oper1[48], g48[32]);
AN2 GA48_33(oper2[33], oper1[48], g48[33]);
AN2 GA48_34(oper2[34], oper1[48], g48[34]);
AN2 GA48_35(oper2[35], oper1[48], g48[35]);
AN2 GA48_36(oper2[36], oper1[48], g48[36]);
AN2 GA48_37(oper2[37], oper1[48], g48[37]);
AN2 GA48_38(oper2[38], oper1[48], g48[38]);
AN2 GA48_39(oper2[39], oper1[48], g48[39]);
AN2 GA48_40(oper2[40], oper1[48], g48[40]);
AN2 GA48_41(oper2[41], oper1[48], g48[41]);
AN2 GA48_42(oper2[42], oper1[48], g48[42]);
AN2 GA48_43(oper2[43], oper1[48], g48[43]);
AN2 GA48_44(oper2[44], oper1[48], g48[44]);
AN2 GA48_45(oper2[45], oper1[48], g48[45]);
AN2 GA48_46(oper2[46], oper1[48], g48[46]);
AN2 GA48_47(oper2[47], oper1[48], g48[47]);
AN2 GA48_48(oper2[48], oper1[48], g48[48]);
AN2 GA48_49(oper2[49], oper1[48], g48[49]);
AN2 GA48_50(oper2[50], oper1[48], g48[50]);
AN2 GA48_51(oper2[51], oper1[48], g48[51]);
AN2 GA48_52(oper2[52], oper1[48], g48[52]);
AN2 GA48_53(oper2[53], oper1[48], g48[53]);
AN2 GA48_54(oper2[54], oper1[48], g48[54]);
AN2 GA48_55(oper2[55], oper1[48], g48[55]);
AN2 GA48_56(oper2[56], oper1[48], g48[56]);
AN2 GA48_57(oper2[57], oper1[48], g48[57]);
AN2 GA48_58(oper2[58], oper1[48], g48[58]);
AN2 GA48_59(oper2[59], oper1[48], g48[59]);
AN2 GA48_60(oper2[60], oper1[48], g48[60]);
AN2 GA48_61(oper2[61], oper1[48], g48[61]);
AN2 GA48_62(oper2[62], oper1[48], g48[62]);
AN2 GA48_63(oper2[63], oper1[48], g48[63]);
AN2 GA47_8(oper2[8], oper1[47], g47[8]);
AN2 GA47_9(oper2[9], oper1[47], g47[9]);
AN2 GA47_10(oper2[10], oper1[47], g47[10]);
AN2 GA47_11(oper2[11], oper1[47], g47[11]);
AN2 GA47_12(oper2[12], oper1[47], g47[12]);
AN2 GA47_13(oper2[13], oper1[47], g47[13]);
AN2 GA47_14(oper2[14], oper1[47], g47[14]);
AN2 GA47_15(oper2[15], oper1[47], g47[15]);
AN2 GA47_16(oper2[16], oper1[47], g47[16]);
AN2 GA47_17(oper2[17], oper1[47], g47[17]);
AN2 GA47_18(oper2[18], oper1[47], g47[18]);
AN2 GA47_19(oper2[19], oper1[47], g47[19]);
AN2 GA47_20(oper2[20], oper1[47], g47[20]);
AN2 GA47_21(oper2[21], oper1[47], g47[21]);
AN2 GA47_22(oper2[22], oper1[47], g47[22]);
AN2 GA47_23(oper2[23], oper1[47], g47[23]);
AN2 GA47_24(oper2[24], oper1[47], g47[24]);
AN2 GA47_25(oper2[25], oper1[47], g47[25]);
AN2 GA47_26(oper2[26], oper1[47], g47[26]);
AN2 GA47_27(oper2[27], oper1[47], g47[27]);
AN2 GA47_28(oper2[28], oper1[47], g47[28]);
AN2 GA47_29(oper2[29], oper1[47], g47[29]);
AN2 GA47_30(oper2[30], oper1[47], g47[30]);
AN2 GA47_31(oper2[31], oper1[47], g47[31]);
AN2 GA47_32(oper2[32], oper1[47], g47[32]);
AN2 GA47_33(oper2[33], oper1[47], g47[33]);
AN2 GA47_34(oper2[34], oper1[47], g47[34]);
AN2 GA47_35(oper2[35], oper1[47], g47[35]);
AN2 GA47_36(oper2[36], oper1[47], g47[36]);
AN2 GA47_37(oper2[37], oper1[47], g47[37]);
AN2 GA47_38(oper2[38], oper1[47], g47[38]);
AN2 GA47_39(oper2[39], oper1[47], g47[39]);
AN2 GA47_40(oper2[40], oper1[47], g47[40]);
AN2 GA47_41(oper2[41], oper1[47], g47[41]);
AN2 GA47_42(oper2[42], oper1[47], g47[42]);
AN2 GA47_43(oper2[43], oper1[47], g47[43]);
AN2 GA47_44(oper2[44], oper1[47], g47[44]);
AN2 GA47_45(oper2[45], oper1[47], g47[45]);
AN2 GA47_46(oper2[46], oper1[47], g47[46]);
AN2 GA47_47(oper2[47], oper1[47], g47[47]);
AN2 GA47_48(oper2[48], oper1[47], g47[48]);
AN2 GA47_49(oper2[49], oper1[47], g47[49]);
AN2 GA47_50(oper2[50], oper1[47], g47[50]);
AN2 GA47_51(oper2[51], oper1[47], g47[51]);
AN2 GA47_52(oper2[52], oper1[47], g47[52]);
AN2 GA47_53(oper2[53], oper1[47], g47[53]);
AN2 GA47_54(oper2[54], oper1[47], g47[54]);
AN2 GA47_55(oper2[55], oper1[47], g47[55]);
AN2 GA47_56(oper2[56], oper1[47], g47[56]);
AN2 GA47_57(oper2[57], oper1[47], g47[57]);
AN2 GA47_58(oper2[58], oper1[47], g47[58]);
AN2 GA47_59(oper2[59], oper1[47], g47[59]);
AN2 GA47_60(oper2[60], oper1[47], g47[60]);
AN2 GA47_61(oper2[61], oper1[47], g47[61]);
AN2 GA47_62(oper2[62], oper1[47], g47[62]);
AN2 GA47_63(oper2[63], oper1[47], g47[63]);
AN2 GA46_8(oper2[8], oper1[46], g46[8]);
AN2 GA46_9(oper2[9], oper1[46], g46[9]);
AN2 GA46_10(oper2[10], oper1[46], g46[10]);
AN2 GA46_11(oper2[11], oper1[46], g46[11]);
AN2 GA46_12(oper2[12], oper1[46], g46[12]);
AN2 GA46_13(oper2[13], oper1[46], g46[13]);
AN2 GA46_14(oper2[14], oper1[46], g46[14]);
AN2 GA46_15(oper2[15], oper1[46], g46[15]);
AN2 GA46_16(oper2[16], oper1[46], g46[16]);
AN2 GA46_17(oper2[17], oper1[46], g46[17]);
AN2 GA46_18(oper2[18], oper1[46], g46[18]);
AN2 GA46_19(oper2[19], oper1[46], g46[19]);
AN2 GA46_20(oper2[20], oper1[46], g46[20]);
AN2 GA46_21(oper2[21], oper1[46], g46[21]);
AN2 GA46_22(oper2[22], oper1[46], g46[22]);
AN2 GA46_23(oper2[23], oper1[46], g46[23]);
AN2 GA46_24(oper2[24], oper1[46], g46[24]);
AN2 GA46_25(oper2[25], oper1[46], g46[25]);
AN2 GA46_26(oper2[26], oper1[46], g46[26]);
AN2 GA46_27(oper2[27], oper1[46], g46[27]);
AN2 GA46_28(oper2[28], oper1[46], g46[28]);
AN2 GA46_29(oper2[29], oper1[46], g46[29]);
AN2 GA46_30(oper2[30], oper1[46], g46[30]);
AN2 GA46_31(oper2[31], oper1[46], g46[31]);
AN2 GA46_32(oper2[32], oper1[46], g46[32]);
AN2 GA46_33(oper2[33], oper1[46], g46[33]);
AN2 GA46_34(oper2[34], oper1[46], g46[34]);
AN2 GA46_35(oper2[35], oper1[46], g46[35]);
AN2 GA46_36(oper2[36], oper1[46], g46[36]);
AN2 GA46_37(oper2[37], oper1[46], g46[37]);
AN2 GA46_38(oper2[38], oper1[46], g46[38]);
AN2 GA46_39(oper2[39], oper1[46], g46[39]);
AN2 GA46_40(oper2[40], oper1[46], g46[40]);
AN2 GA46_41(oper2[41], oper1[46], g46[41]);
AN2 GA46_42(oper2[42], oper1[46], g46[42]);
AN2 GA46_43(oper2[43], oper1[46], g46[43]);
AN2 GA46_44(oper2[44], oper1[46], g46[44]);
AN2 GA46_45(oper2[45], oper1[46], g46[45]);
AN2 GA46_46(oper2[46], oper1[46], g46[46]);
AN2 GA46_47(oper2[47], oper1[46], g46[47]);
AN2 GA46_48(oper2[48], oper1[46], g46[48]);
AN2 GA46_49(oper2[49], oper1[46], g46[49]);
AN2 GA46_50(oper2[50], oper1[46], g46[50]);
AN2 GA46_51(oper2[51], oper1[46], g46[51]);
AN2 GA46_52(oper2[52], oper1[46], g46[52]);
AN2 GA46_53(oper2[53], oper1[46], g46[53]);
AN2 GA46_54(oper2[54], oper1[46], g46[54]);
AN2 GA46_55(oper2[55], oper1[46], g46[55]);
AN2 GA46_56(oper2[56], oper1[46], g46[56]);
AN2 GA46_57(oper2[57], oper1[46], g46[57]);
AN2 GA46_58(oper2[58], oper1[46], g46[58]);
AN2 GA46_59(oper2[59], oper1[46], g46[59]);
AN2 GA46_60(oper2[60], oper1[46], g46[60]);
AN2 GA46_61(oper2[61], oper1[46], g46[61]);
AN2 GA46_62(oper2[62], oper1[46], g46[62]);
AN2 GA46_63(oper2[63], oper1[46], g46[63]);
AN2 GA45_8(oper2[8], oper1[45], g45[8]);
AN2 GA45_9(oper2[9], oper1[45], g45[9]);
AN2 GA45_10(oper2[10], oper1[45], g45[10]);
AN2 GA45_11(oper2[11], oper1[45], g45[11]);
AN2 GA45_12(oper2[12], oper1[45], g45[12]);
AN2 GA45_13(oper2[13], oper1[45], g45[13]);
AN2 GA45_14(oper2[14], oper1[45], g45[14]);
AN2 GA45_15(oper2[15], oper1[45], g45[15]);
AN2 GA45_16(oper2[16], oper1[45], g45[16]);
AN2 GA45_17(oper2[17], oper1[45], g45[17]);
AN2 GA45_18(oper2[18], oper1[45], g45[18]);
AN2 GA45_19(oper2[19], oper1[45], g45[19]);
AN2 GA45_20(oper2[20], oper1[45], g45[20]);
AN2 GA45_21(oper2[21], oper1[45], g45[21]);
AN2 GA45_22(oper2[22], oper1[45], g45[22]);
AN2 GA45_23(oper2[23], oper1[45], g45[23]);
AN2 GA45_24(oper2[24], oper1[45], g45[24]);
AN2 GA45_25(oper2[25], oper1[45], g45[25]);
AN2 GA45_26(oper2[26], oper1[45], g45[26]);
AN2 GA45_27(oper2[27], oper1[45], g45[27]);
AN2 GA45_28(oper2[28], oper1[45], g45[28]);
AN2 GA45_29(oper2[29], oper1[45], g45[29]);
AN2 GA45_30(oper2[30], oper1[45], g45[30]);
AN2 GA45_31(oper2[31], oper1[45], g45[31]);
AN2 GA45_32(oper2[32], oper1[45], g45[32]);
AN2 GA45_33(oper2[33], oper1[45], g45[33]);
AN2 GA45_34(oper2[34], oper1[45], g45[34]);
AN2 GA45_35(oper2[35], oper1[45], g45[35]);
AN2 GA45_36(oper2[36], oper1[45], g45[36]);
AN2 GA45_37(oper2[37], oper1[45], g45[37]);
AN2 GA45_38(oper2[38], oper1[45], g45[38]);
AN2 GA45_39(oper2[39], oper1[45], g45[39]);
AN2 GA45_40(oper2[40], oper1[45], g45[40]);
AN2 GA45_41(oper2[41], oper1[45], g45[41]);
AN2 GA45_42(oper2[42], oper1[45], g45[42]);
AN2 GA45_43(oper2[43], oper1[45], g45[43]);
AN2 GA45_44(oper2[44], oper1[45], g45[44]);
AN2 GA45_45(oper2[45], oper1[45], g45[45]);
AN2 GA45_46(oper2[46], oper1[45], g45[46]);
AN2 GA45_47(oper2[47], oper1[45], g45[47]);
AN2 GA45_48(oper2[48], oper1[45], g45[48]);
AN2 GA45_49(oper2[49], oper1[45], g45[49]);
AN2 GA45_50(oper2[50], oper1[45], g45[50]);
AN2 GA45_51(oper2[51], oper1[45], g45[51]);
AN2 GA45_52(oper2[52], oper1[45], g45[52]);
AN2 GA45_53(oper2[53], oper1[45], g45[53]);
AN2 GA45_54(oper2[54], oper1[45], g45[54]);
AN2 GA45_55(oper2[55], oper1[45], g45[55]);
AN2 GA45_56(oper2[56], oper1[45], g45[56]);
AN2 GA45_57(oper2[57], oper1[45], g45[57]);
AN2 GA45_58(oper2[58], oper1[45], g45[58]);
AN2 GA45_59(oper2[59], oper1[45], g45[59]);
AN2 GA45_60(oper2[60], oper1[45], g45[60]);
AN2 GA45_61(oper2[61], oper1[45], g45[61]);
AN2 GA45_62(oper2[62], oper1[45], g45[62]);
AN2 GA45_63(oper2[63], oper1[45], g45[63]);
AN2 GA44_8(oper2[8], oper1[44], g44[8]);
AN2 GA44_9(oper2[9], oper1[44], g44[9]);
AN2 GA44_10(oper2[10], oper1[44], g44[10]);
AN2 GA44_11(oper2[11], oper1[44], g44[11]);
AN2 GA44_12(oper2[12], oper1[44], g44[12]);
AN2 GA44_13(oper2[13], oper1[44], g44[13]);
AN2 GA44_14(oper2[14], oper1[44], g44[14]);
AN2 GA44_15(oper2[15], oper1[44], g44[15]);
AN2 GA44_16(oper2[16], oper1[44], g44[16]);
AN2 GA44_17(oper2[17], oper1[44], g44[17]);
AN2 GA44_18(oper2[18], oper1[44], g44[18]);
AN2 GA44_19(oper2[19], oper1[44], g44[19]);
AN2 GA44_20(oper2[20], oper1[44], g44[20]);
AN2 GA44_21(oper2[21], oper1[44], g44[21]);
AN2 GA44_22(oper2[22], oper1[44], g44[22]);
AN2 GA44_23(oper2[23], oper1[44], g44[23]);
AN2 GA44_24(oper2[24], oper1[44], g44[24]);
AN2 GA44_25(oper2[25], oper1[44], g44[25]);
AN2 GA44_26(oper2[26], oper1[44], g44[26]);
AN2 GA44_27(oper2[27], oper1[44], g44[27]);
AN2 GA44_28(oper2[28], oper1[44], g44[28]);
AN2 GA44_29(oper2[29], oper1[44], g44[29]);
AN2 GA44_30(oper2[30], oper1[44], g44[30]);
AN2 GA44_31(oper2[31], oper1[44], g44[31]);
AN2 GA44_32(oper2[32], oper1[44], g44[32]);
AN2 GA44_33(oper2[33], oper1[44], g44[33]);
AN2 GA44_34(oper2[34], oper1[44], g44[34]);
AN2 GA44_35(oper2[35], oper1[44], g44[35]);
AN2 GA44_36(oper2[36], oper1[44], g44[36]);
AN2 GA44_37(oper2[37], oper1[44], g44[37]);
AN2 GA44_38(oper2[38], oper1[44], g44[38]);
AN2 GA44_39(oper2[39], oper1[44], g44[39]);
AN2 GA44_40(oper2[40], oper1[44], g44[40]);
AN2 GA44_41(oper2[41], oper1[44], g44[41]);
AN2 GA44_42(oper2[42], oper1[44], g44[42]);
AN2 GA44_43(oper2[43], oper1[44], g44[43]);
AN2 GA44_44(oper2[44], oper1[44], g44[44]);
AN2 GA44_45(oper2[45], oper1[44], g44[45]);
AN2 GA44_46(oper2[46], oper1[44], g44[46]);
AN2 GA44_47(oper2[47], oper1[44], g44[47]);
AN2 GA44_48(oper2[48], oper1[44], g44[48]);
AN2 GA44_49(oper2[49], oper1[44], g44[49]);
AN2 GA44_50(oper2[50], oper1[44], g44[50]);
AN2 GA44_51(oper2[51], oper1[44], g44[51]);
AN2 GA44_52(oper2[52], oper1[44], g44[52]);
AN2 GA44_53(oper2[53], oper1[44], g44[53]);
AN2 GA44_54(oper2[54], oper1[44], g44[54]);
AN2 GA44_55(oper2[55], oper1[44], g44[55]);
AN2 GA44_56(oper2[56], oper1[44], g44[56]);
AN2 GA44_57(oper2[57], oper1[44], g44[57]);
AN2 GA44_58(oper2[58], oper1[44], g44[58]);
AN2 GA44_59(oper2[59], oper1[44], g44[59]);
AN2 GA44_60(oper2[60], oper1[44], g44[60]);
AN2 GA44_61(oper2[61], oper1[44], g44[61]);
AN2 GA44_62(oper2[62], oper1[44], g44[62]);
AN2 GA44_63(oper2[63], oper1[44], g44[63]);
AN2 GA43_8(oper2[8], oper1[43], g43[8]);
AN2 GA43_9(oper2[9], oper1[43], g43[9]);
AN2 GA43_10(oper2[10], oper1[43], g43[10]);
AN2 GA43_11(oper2[11], oper1[43], g43[11]);
AN2 GA43_12(oper2[12], oper1[43], g43[12]);
AN2 GA43_13(oper2[13], oper1[43], g43[13]);
AN2 GA43_14(oper2[14], oper1[43], g43[14]);
AN2 GA43_15(oper2[15], oper1[43], g43[15]);
AN2 GA43_16(oper2[16], oper1[43], g43[16]);
AN2 GA43_17(oper2[17], oper1[43], g43[17]);
AN2 GA43_18(oper2[18], oper1[43], g43[18]);
AN2 GA43_19(oper2[19], oper1[43], g43[19]);
AN2 GA43_20(oper2[20], oper1[43], g43[20]);
AN2 GA43_21(oper2[21], oper1[43], g43[21]);
AN2 GA43_22(oper2[22], oper1[43], g43[22]);
AN2 GA43_23(oper2[23], oper1[43], g43[23]);
AN2 GA43_24(oper2[24], oper1[43], g43[24]);
AN2 GA43_25(oper2[25], oper1[43], g43[25]);
AN2 GA43_26(oper2[26], oper1[43], g43[26]);
AN2 GA43_27(oper2[27], oper1[43], g43[27]);
AN2 GA43_28(oper2[28], oper1[43], g43[28]);
AN2 GA43_29(oper2[29], oper1[43], g43[29]);
AN2 GA43_30(oper2[30], oper1[43], g43[30]);
AN2 GA43_31(oper2[31], oper1[43], g43[31]);
AN2 GA43_32(oper2[32], oper1[43], g43[32]);
AN2 GA43_33(oper2[33], oper1[43], g43[33]);
AN2 GA43_34(oper2[34], oper1[43], g43[34]);
AN2 GA43_35(oper2[35], oper1[43], g43[35]);
AN2 GA43_36(oper2[36], oper1[43], g43[36]);
AN2 GA43_37(oper2[37], oper1[43], g43[37]);
AN2 GA43_38(oper2[38], oper1[43], g43[38]);
AN2 GA43_39(oper2[39], oper1[43], g43[39]);
AN2 GA43_40(oper2[40], oper1[43], g43[40]);
AN2 GA43_41(oper2[41], oper1[43], g43[41]);
AN2 GA43_42(oper2[42], oper1[43], g43[42]);
AN2 GA43_43(oper2[43], oper1[43], g43[43]);
AN2 GA43_44(oper2[44], oper1[43], g43[44]);
AN2 GA43_45(oper2[45], oper1[43], g43[45]);
AN2 GA43_46(oper2[46], oper1[43], g43[46]);
AN2 GA43_47(oper2[47], oper1[43], g43[47]);
AN2 GA43_48(oper2[48], oper1[43], g43[48]);
AN2 GA43_49(oper2[49], oper1[43], g43[49]);
AN2 GA43_50(oper2[50], oper1[43], g43[50]);
AN2 GA43_51(oper2[51], oper1[43], g43[51]);
AN2 GA43_52(oper2[52], oper1[43], g43[52]);
AN2 GA43_53(oper2[53], oper1[43], g43[53]);
AN2 GA43_54(oper2[54], oper1[43], g43[54]);
AN2 GA43_55(oper2[55], oper1[43], g43[55]);
AN2 GA43_56(oper2[56], oper1[43], g43[56]);
AN2 GA43_57(oper2[57], oper1[43], g43[57]);
AN2 GA43_58(oper2[58], oper1[43], g43[58]);
AN2 GA43_59(oper2[59], oper1[43], g43[59]);
AN2 GA43_60(oper2[60], oper1[43], g43[60]);
AN2 GA43_61(oper2[61], oper1[43], g43[61]);
AN2 GA43_62(oper2[62], oper1[43], g43[62]);
AN2 GA43_63(oper2[63], oper1[43], g43[63]);
AN2 GA42_8(oper2[8], oper1[42], g42[8]);
AN2 GA42_9(oper2[9], oper1[42], g42[9]);
AN2 GA42_10(oper2[10], oper1[42], g42[10]);
AN2 GA42_11(oper2[11], oper1[42], g42[11]);
AN2 GA42_12(oper2[12], oper1[42], g42[12]);
AN2 GA42_13(oper2[13], oper1[42], g42[13]);
AN2 GA42_14(oper2[14], oper1[42], g42[14]);
AN2 GA42_15(oper2[15], oper1[42], g42[15]);
AN2 GA42_16(oper2[16], oper1[42], g42[16]);
AN2 GA42_17(oper2[17], oper1[42], g42[17]);
AN2 GA42_18(oper2[18], oper1[42], g42[18]);
AN2 GA42_19(oper2[19], oper1[42], g42[19]);
AN2 GA42_20(oper2[20], oper1[42], g42[20]);
AN2 GA42_21(oper2[21], oper1[42], g42[21]);
AN2 GA42_22(oper2[22], oper1[42], g42[22]);
AN2 GA42_23(oper2[23], oper1[42], g42[23]);
AN2 GA42_24(oper2[24], oper1[42], g42[24]);
AN2 GA42_25(oper2[25], oper1[42], g42[25]);
AN2 GA42_26(oper2[26], oper1[42], g42[26]);
AN2 GA42_27(oper2[27], oper1[42], g42[27]);
AN2 GA42_28(oper2[28], oper1[42], g42[28]);
AN2 GA42_29(oper2[29], oper1[42], g42[29]);
AN2 GA42_30(oper2[30], oper1[42], g42[30]);
AN2 GA42_31(oper2[31], oper1[42], g42[31]);
AN2 GA42_32(oper2[32], oper1[42], g42[32]);
AN2 GA42_33(oper2[33], oper1[42], g42[33]);
AN2 GA42_34(oper2[34], oper1[42], g42[34]);
AN2 GA42_35(oper2[35], oper1[42], g42[35]);
AN2 GA42_36(oper2[36], oper1[42], g42[36]);
AN2 GA42_37(oper2[37], oper1[42], g42[37]);
AN2 GA42_38(oper2[38], oper1[42], g42[38]);
AN2 GA42_39(oper2[39], oper1[42], g42[39]);
AN2 GA42_40(oper2[40], oper1[42], g42[40]);
AN2 GA42_41(oper2[41], oper1[42], g42[41]);
AN2 GA42_42(oper2[42], oper1[42], g42[42]);
AN2 GA42_43(oper2[43], oper1[42], g42[43]);
AN2 GA42_44(oper2[44], oper1[42], g42[44]);
AN2 GA42_45(oper2[45], oper1[42], g42[45]);
AN2 GA42_46(oper2[46], oper1[42], g42[46]);
AN2 GA42_47(oper2[47], oper1[42], g42[47]);
AN2 GA42_48(oper2[48], oper1[42], g42[48]);
AN2 GA42_49(oper2[49], oper1[42], g42[49]);
AN2 GA42_50(oper2[50], oper1[42], g42[50]);
AN2 GA42_51(oper2[51], oper1[42], g42[51]);
AN2 GA42_52(oper2[52], oper1[42], g42[52]);
AN2 GA42_53(oper2[53], oper1[42], g42[53]);
AN2 GA42_54(oper2[54], oper1[42], g42[54]);
AN2 GA42_55(oper2[55], oper1[42], g42[55]);
AN2 GA42_56(oper2[56], oper1[42], g42[56]);
AN2 GA42_57(oper2[57], oper1[42], g42[57]);
AN2 GA42_58(oper2[58], oper1[42], g42[58]);
AN2 GA42_59(oper2[59], oper1[42], g42[59]);
AN2 GA42_60(oper2[60], oper1[42], g42[60]);
AN2 GA42_61(oper2[61], oper1[42], g42[61]);
AN2 GA42_62(oper2[62], oper1[42], g42[62]);
AN2 GA42_63(oper2[63], oper1[42], g42[63]);
AN2 GA41_8(oper2[8], oper1[41], g41[8]);
AN2 GA41_9(oper2[9], oper1[41], g41[9]);
AN2 GA41_10(oper2[10], oper1[41], g41[10]);
AN2 GA41_11(oper2[11], oper1[41], g41[11]);
AN2 GA41_12(oper2[12], oper1[41], g41[12]);
AN2 GA41_13(oper2[13], oper1[41], g41[13]);
AN2 GA41_14(oper2[14], oper1[41], g41[14]);
AN2 GA41_15(oper2[15], oper1[41], g41[15]);
AN2 GA41_16(oper2[16], oper1[41], g41[16]);
AN2 GA41_17(oper2[17], oper1[41], g41[17]);
AN2 GA41_18(oper2[18], oper1[41], g41[18]);
AN2 GA41_19(oper2[19], oper1[41], g41[19]);
AN2 GA41_20(oper2[20], oper1[41], g41[20]);
AN2 GA41_21(oper2[21], oper1[41], g41[21]);
AN2 GA41_22(oper2[22], oper1[41], g41[22]);
AN2 GA41_23(oper2[23], oper1[41], g41[23]);
AN2 GA41_24(oper2[24], oper1[41], g41[24]);
AN2 GA41_25(oper2[25], oper1[41], g41[25]);
AN2 GA41_26(oper2[26], oper1[41], g41[26]);
AN2 GA41_27(oper2[27], oper1[41], g41[27]);
AN2 GA41_28(oper2[28], oper1[41], g41[28]);
AN2 GA41_29(oper2[29], oper1[41], g41[29]);
AN2 GA41_30(oper2[30], oper1[41], g41[30]);
AN2 GA41_31(oper2[31], oper1[41], g41[31]);
AN2 GA41_32(oper2[32], oper1[41], g41[32]);
AN2 GA41_33(oper2[33], oper1[41], g41[33]);
AN2 GA41_34(oper2[34], oper1[41], g41[34]);
AN2 GA41_35(oper2[35], oper1[41], g41[35]);
AN2 GA41_36(oper2[36], oper1[41], g41[36]);
AN2 GA41_37(oper2[37], oper1[41], g41[37]);
AN2 GA41_38(oper2[38], oper1[41], g41[38]);
AN2 GA41_39(oper2[39], oper1[41], g41[39]);
AN2 GA41_40(oper2[40], oper1[41], g41[40]);
AN2 GA41_41(oper2[41], oper1[41], g41[41]);
AN2 GA41_42(oper2[42], oper1[41], g41[42]);
AN2 GA41_43(oper2[43], oper1[41], g41[43]);
AN2 GA41_44(oper2[44], oper1[41], g41[44]);
AN2 GA41_45(oper2[45], oper1[41], g41[45]);
AN2 GA41_46(oper2[46], oper1[41], g41[46]);
AN2 GA41_47(oper2[47], oper1[41], g41[47]);
AN2 GA41_48(oper2[48], oper1[41], g41[48]);
AN2 GA41_49(oper2[49], oper1[41], g41[49]);
AN2 GA41_50(oper2[50], oper1[41], g41[50]);
AN2 GA41_51(oper2[51], oper1[41], g41[51]);
AN2 GA41_52(oper2[52], oper1[41], g41[52]);
AN2 GA41_53(oper2[53], oper1[41], g41[53]);
AN2 GA41_54(oper2[54], oper1[41], g41[54]);
AN2 GA41_55(oper2[55], oper1[41], g41[55]);
AN2 GA41_56(oper2[56], oper1[41], g41[56]);
AN2 GA41_57(oper2[57], oper1[41], g41[57]);
AN2 GA41_58(oper2[58], oper1[41], g41[58]);
AN2 GA41_59(oper2[59], oper1[41], g41[59]);
AN2 GA41_60(oper2[60], oper1[41], g41[60]);
AN2 GA41_61(oper2[61], oper1[41], g41[61]);
AN2 GA41_62(oper2[62], oper1[41], g41[62]);
AN2 GA41_63(oper2[63], oper1[41], g41[63]);
AN2 GA40_8(oper2[8], oper1[40], g40[8]);
AN2 GA40_9(oper2[9], oper1[40], g40[9]);
AN2 GA40_10(oper2[10], oper1[40], g40[10]);
AN2 GA40_11(oper2[11], oper1[40], g40[11]);
AN2 GA40_12(oper2[12], oper1[40], g40[12]);
AN2 GA40_13(oper2[13], oper1[40], g40[13]);
AN2 GA40_14(oper2[14], oper1[40], g40[14]);
AN2 GA40_15(oper2[15], oper1[40], g40[15]);
AN2 GA40_16(oper2[16], oper1[40], g40[16]);
AN2 GA40_17(oper2[17], oper1[40], g40[17]);
AN2 GA40_18(oper2[18], oper1[40], g40[18]);
AN2 GA40_19(oper2[19], oper1[40], g40[19]);
AN2 GA40_20(oper2[20], oper1[40], g40[20]);
AN2 GA40_21(oper2[21], oper1[40], g40[21]);
AN2 GA40_22(oper2[22], oper1[40], g40[22]);
AN2 GA40_23(oper2[23], oper1[40], g40[23]);
AN2 GA40_24(oper2[24], oper1[40], g40[24]);
AN2 GA40_25(oper2[25], oper1[40], g40[25]);
AN2 GA40_26(oper2[26], oper1[40], g40[26]);
AN2 GA40_27(oper2[27], oper1[40], g40[27]);
AN2 GA40_28(oper2[28], oper1[40], g40[28]);
AN2 GA40_29(oper2[29], oper1[40], g40[29]);
AN2 GA40_30(oper2[30], oper1[40], g40[30]);
AN2 GA40_31(oper2[31], oper1[40], g40[31]);
AN2 GA40_32(oper2[32], oper1[40], g40[32]);
AN2 GA40_33(oper2[33], oper1[40], g40[33]);
AN2 GA40_34(oper2[34], oper1[40], g40[34]);
AN2 GA40_35(oper2[35], oper1[40], g40[35]);
AN2 GA40_36(oper2[36], oper1[40], g40[36]);
AN2 GA40_37(oper2[37], oper1[40], g40[37]);
AN2 GA40_38(oper2[38], oper1[40], g40[38]);
AN2 GA40_39(oper2[39], oper1[40], g40[39]);
AN2 GA40_40(oper2[40], oper1[40], g40[40]);
AN2 GA40_41(oper2[41], oper1[40], g40[41]);
AN2 GA40_42(oper2[42], oper1[40], g40[42]);
AN2 GA40_43(oper2[43], oper1[40], g40[43]);
AN2 GA40_44(oper2[44], oper1[40], g40[44]);
AN2 GA40_45(oper2[45], oper1[40], g40[45]);
AN2 GA40_46(oper2[46], oper1[40], g40[46]);
AN2 GA40_47(oper2[47], oper1[40], g40[47]);
AN2 GA40_48(oper2[48], oper1[40], g40[48]);
AN2 GA40_49(oper2[49], oper1[40], g40[49]);
AN2 GA40_50(oper2[50], oper1[40], g40[50]);
AN2 GA40_51(oper2[51], oper1[40], g40[51]);
AN2 GA40_52(oper2[52], oper1[40], g40[52]);
AN2 GA40_53(oper2[53], oper1[40], g40[53]);
AN2 GA40_54(oper2[54], oper1[40], g40[54]);
AN2 GA40_55(oper2[55], oper1[40], g40[55]);
AN2 GA40_56(oper2[56], oper1[40], g40[56]);
AN2 GA40_57(oper2[57], oper1[40], g40[57]);
AN2 GA40_58(oper2[58], oper1[40], g40[58]);
AN2 GA40_59(oper2[59], oper1[40], g40[59]);
AN2 GA40_60(oper2[60], oper1[40], g40[60]);
AN2 GA40_61(oper2[61], oper1[40], g40[61]);
AN2 GA40_62(oper2[62], oper1[40], g40[62]);
AN2 GA40_63(oper2[63], oper1[40], g40[63]);
AN2 GA39_8(oper2[8], oper1[39], g39[8]);
AN2 GA39_9(oper2[9], oper1[39], g39[9]);
AN2 GA39_10(oper2[10], oper1[39], g39[10]);
AN2 GA39_11(oper2[11], oper1[39], g39[11]);
AN2 GA39_12(oper2[12], oper1[39], g39[12]);
AN2 GA39_13(oper2[13], oper1[39], g39[13]);
AN2 GA39_14(oper2[14], oper1[39], g39[14]);
AN2 GA39_15(oper2[15], oper1[39], g39[15]);
AN2 GA39_16(oper2[16], oper1[39], g39[16]);
AN2 GA39_17(oper2[17], oper1[39], g39[17]);
AN2 GA39_18(oper2[18], oper1[39], g39[18]);
AN2 GA39_19(oper2[19], oper1[39], g39[19]);
AN2 GA39_20(oper2[20], oper1[39], g39[20]);
AN2 GA39_21(oper2[21], oper1[39], g39[21]);
AN2 GA39_22(oper2[22], oper1[39], g39[22]);
AN2 GA39_23(oper2[23], oper1[39], g39[23]);
AN2 GA39_24(oper2[24], oper1[39], g39[24]);
AN2 GA39_25(oper2[25], oper1[39], g39[25]);
AN2 GA39_26(oper2[26], oper1[39], g39[26]);
AN2 GA39_27(oper2[27], oper1[39], g39[27]);
AN2 GA39_28(oper2[28], oper1[39], g39[28]);
AN2 GA39_29(oper2[29], oper1[39], g39[29]);
AN2 GA39_30(oper2[30], oper1[39], g39[30]);
AN2 GA39_31(oper2[31], oper1[39], g39[31]);
AN2 GA39_32(oper2[32], oper1[39], g39[32]);
AN2 GA39_33(oper2[33], oper1[39], g39[33]);
AN2 GA39_34(oper2[34], oper1[39], g39[34]);
AN2 GA39_35(oper2[35], oper1[39], g39[35]);
AN2 GA39_36(oper2[36], oper1[39], g39[36]);
AN2 GA39_37(oper2[37], oper1[39], g39[37]);
AN2 GA39_38(oper2[38], oper1[39], g39[38]);
AN2 GA39_39(oper2[39], oper1[39], g39[39]);
AN2 GA39_40(oper2[40], oper1[39], g39[40]);
AN2 GA39_41(oper2[41], oper1[39], g39[41]);
AN2 GA39_42(oper2[42], oper1[39], g39[42]);
AN2 GA39_43(oper2[43], oper1[39], g39[43]);
AN2 GA39_44(oper2[44], oper1[39], g39[44]);
AN2 GA39_45(oper2[45], oper1[39], g39[45]);
AN2 GA39_46(oper2[46], oper1[39], g39[46]);
AN2 GA39_47(oper2[47], oper1[39], g39[47]);
AN2 GA39_48(oper2[48], oper1[39], g39[48]);
AN2 GA39_49(oper2[49], oper1[39], g39[49]);
AN2 GA39_50(oper2[50], oper1[39], g39[50]);
AN2 GA39_51(oper2[51], oper1[39], g39[51]);
AN2 GA39_52(oper2[52], oper1[39], g39[52]);
AN2 GA39_53(oper2[53], oper1[39], g39[53]);
AN2 GA39_54(oper2[54], oper1[39], g39[54]);
AN2 GA39_55(oper2[55], oper1[39], g39[55]);
AN2 GA39_56(oper2[56], oper1[39], g39[56]);
AN2 GA39_57(oper2[57], oper1[39], g39[57]);
AN2 GA39_58(oper2[58], oper1[39], g39[58]);
AN2 GA39_59(oper2[59], oper1[39], g39[59]);
AN2 GA39_60(oper2[60], oper1[39], g39[60]);
AN2 GA39_61(oper2[61], oper1[39], g39[61]);
AN2 GA39_62(oper2[62], oper1[39], g39[62]);
AN2 GA39_63(oper2[63], oper1[39], g39[63]);
AN2 GA38_8(oper2[8], oper1[38], g38[8]);
AN2 GA38_9(oper2[9], oper1[38], g38[9]);
AN2 GA38_10(oper2[10], oper1[38], g38[10]);
AN2 GA38_11(oper2[11], oper1[38], g38[11]);
AN2 GA38_12(oper2[12], oper1[38], g38[12]);
AN2 GA38_13(oper2[13], oper1[38], g38[13]);
AN2 GA38_14(oper2[14], oper1[38], g38[14]);
AN2 GA38_15(oper2[15], oper1[38], g38[15]);
AN2 GA38_16(oper2[16], oper1[38], g38[16]);
AN2 GA38_17(oper2[17], oper1[38], g38[17]);
AN2 GA38_18(oper2[18], oper1[38], g38[18]);
AN2 GA38_19(oper2[19], oper1[38], g38[19]);
AN2 GA38_20(oper2[20], oper1[38], g38[20]);
AN2 GA38_21(oper2[21], oper1[38], g38[21]);
AN2 GA38_22(oper2[22], oper1[38], g38[22]);
AN2 GA38_23(oper2[23], oper1[38], g38[23]);
AN2 GA38_24(oper2[24], oper1[38], g38[24]);
AN2 GA38_25(oper2[25], oper1[38], g38[25]);
AN2 GA38_26(oper2[26], oper1[38], g38[26]);
AN2 GA38_27(oper2[27], oper1[38], g38[27]);
AN2 GA38_28(oper2[28], oper1[38], g38[28]);
AN2 GA38_29(oper2[29], oper1[38], g38[29]);
AN2 GA38_30(oper2[30], oper1[38], g38[30]);
AN2 GA38_31(oper2[31], oper1[38], g38[31]);
AN2 GA38_32(oper2[32], oper1[38], g38[32]);
AN2 GA38_33(oper2[33], oper1[38], g38[33]);
AN2 GA38_34(oper2[34], oper1[38], g38[34]);
AN2 GA38_35(oper2[35], oper1[38], g38[35]);
AN2 GA38_36(oper2[36], oper1[38], g38[36]);
AN2 GA38_37(oper2[37], oper1[38], g38[37]);
AN2 GA38_38(oper2[38], oper1[38], g38[38]);
AN2 GA38_39(oper2[39], oper1[38], g38[39]);
AN2 GA38_40(oper2[40], oper1[38], g38[40]);
AN2 GA38_41(oper2[41], oper1[38], g38[41]);
AN2 GA38_42(oper2[42], oper1[38], g38[42]);
AN2 GA38_43(oper2[43], oper1[38], g38[43]);
AN2 GA38_44(oper2[44], oper1[38], g38[44]);
AN2 GA38_45(oper2[45], oper1[38], g38[45]);
AN2 GA38_46(oper2[46], oper1[38], g38[46]);
AN2 GA38_47(oper2[47], oper1[38], g38[47]);
AN2 GA38_48(oper2[48], oper1[38], g38[48]);
AN2 GA38_49(oper2[49], oper1[38], g38[49]);
AN2 GA38_50(oper2[50], oper1[38], g38[50]);
AN2 GA38_51(oper2[51], oper1[38], g38[51]);
AN2 GA38_52(oper2[52], oper1[38], g38[52]);
AN2 GA38_53(oper2[53], oper1[38], g38[53]);
AN2 GA38_54(oper2[54], oper1[38], g38[54]);
AN2 GA38_55(oper2[55], oper1[38], g38[55]);
AN2 GA38_56(oper2[56], oper1[38], g38[56]);
AN2 GA38_57(oper2[57], oper1[38], g38[57]);
AN2 GA38_58(oper2[58], oper1[38], g38[58]);
AN2 GA38_59(oper2[59], oper1[38], g38[59]);
AN2 GA38_60(oper2[60], oper1[38], g38[60]);
AN2 GA38_61(oper2[61], oper1[38], g38[61]);
AN2 GA38_62(oper2[62], oper1[38], g38[62]);
AN2 GA38_63(oper2[63], oper1[38], g38[63]);
AN2 GA37_8(oper2[8], oper1[37], g37[8]);
AN2 GA37_9(oper2[9], oper1[37], g37[9]);
AN2 GA37_10(oper2[10], oper1[37], g37[10]);
AN2 GA37_11(oper2[11], oper1[37], g37[11]);
AN2 GA37_12(oper2[12], oper1[37], g37[12]);
AN2 GA37_13(oper2[13], oper1[37], g37[13]);
AN2 GA37_14(oper2[14], oper1[37], g37[14]);
AN2 GA37_15(oper2[15], oper1[37], g37[15]);
AN2 GA37_16(oper2[16], oper1[37], g37[16]);
AN2 GA37_17(oper2[17], oper1[37], g37[17]);
AN2 GA37_18(oper2[18], oper1[37], g37[18]);
AN2 GA37_19(oper2[19], oper1[37], g37[19]);
AN2 GA37_20(oper2[20], oper1[37], g37[20]);
AN2 GA37_21(oper2[21], oper1[37], g37[21]);
AN2 GA37_22(oper2[22], oper1[37], g37[22]);
AN2 GA37_23(oper2[23], oper1[37], g37[23]);
AN2 GA37_24(oper2[24], oper1[37], g37[24]);
AN2 GA37_25(oper2[25], oper1[37], g37[25]);
AN2 GA37_26(oper2[26], oper1[37], g37[26]);
AN2 GA37_27(oper2[27], oper1[37], g37[27]);
AN2 GA37_28(oper2[28], oper1[37], g37[28]);
AN2 GA37_29(oper2[29], oper1[37], g37[29]);
AN2 GA37_30(oper2[30], oper1[37], g37[30]);
AN2 GA37_31(oper2[31], oper1[37], g37[31]);
AN2 GA37_32(oper2[32], oper1[37], g37[32]);
AN2 GA37_33(oper2[33], oper1[37], g37[33]);
AN2 GA37_34(oper2[34], oper1[37], g37[34]);
AN2 GA37_35(oper2[35], oper1[37], g37[35]);
AN2 GA37_36(oper2[36], oper1[37], g37[36]);
AN2 GA37_37(oper2[37], oper1[37], g37[37]);
AN2 GA37_38(oper2[38], oper1[37], g37[38]);
AN2 GA37_39(oper2[39], oper1[37], g37[39]);
AN2 GA37_40(oper2[40], oper1[37], g37[40]);
AN2 GA37_41(oper2[41], oper1[37], g37[41]);
AN2 GA37_42(oper2[42], oper1[37], g37[42]);
AN2 GA37_43(oper2[43], oper1[37], g37[43]);
AN2 GA37_44(oper2[44], oper1[37], g37[44]);
AN2 GA37_45(oper2[45], oper1[37], g37[45]);
AN2 GA37_46(oper2[46], oper1[37], g37[46]);
AN2 GA37_47(oper2[47], oper1[37], g37[47]);
AN2 GA37_48(oper2[48], oper1[37], g37[48]);
AN2 GA37_49(oper2[49], oper1[37], g37[49]);
AN2 GA37_50(oper2[50], oper1[37], g37[50]);
AN2 GA37_51(oper2[51], oper1[37], g37[51]);
AN2 GA37_52(oper2[52], oper1[37], g37[52]);
AN2 GA37_53(oper2[53], oper1[37], g37[53]);
AN2 GA37_54(oper2[54], oper1[37], g37[54]);
AN2 GA37_55(oper2[55], oper1[37], g37[55]);
AN2 GA37_56(oper2[56], oper1[37], g37[56]);
AN2 GA37_57(oper2[57], oper1[37], g37[57]);
AN2 GA37_58(oper2[58], oper1[37], g37[58]);
AN2 GA37_59(oper2[59], oper1[37], g37[59]);
AN2 GA37_60(oper2[60], oper1[37], g37[60]);
AN2 GA37_61(oper2[61], oper1[37], g37[61]);
AN2 GA37_62(oper2[62], oper1[37], g37[62]);
AN2 GA37_63(oper2[63], oper1[37], g37[63]);
AN2 GA36_8(oper2[8], oper1[36], g36[8]);
AN2 GA36_9(oper2[9], oper1[36], g36[9]);
AN2 GA36_10(oper2[10], oper1[36], g36[10]);
AN2 GA36_11(oper2[11], oper1[36], g36[11]);
AN2 GA36_12(oper2[12], oper1[36], g36[12]);
AN2 GA36_13(oper2[13], oper1[36], g36[13]);
AN2 GA36_14(oper2[14], oper1[36], g36[14]);
AN2 GA36_15(oper2[15], oper1[36], g36[15]);
AN2 GA36_16(oper2[16], oper1[36], g36[16]);
AN2 GA36_17(oper2[17], oper1[36], g36[17]);
AN2 GA36_18(oper2[18], oper1[36], g36[18]);
AN2 GA36_19(oper2[19], oper1[36], g36[19]);
AN2 GA36_20(oper2[20], oper1[36], g36[20]);
AN2 GA36_21(oper2[21], oper1[36], g36[21]);
AN2 GA36_22(oper2[22], oper1[36], g36[22]);
AN2 GA36_23(oper2[23], oper1[36], g36[23]);
AN2 GA36_24(oper2[24], oper1[36], g36[24]);
AN2 GA36_25(oper2[25], oper1[36], g36[25]);
AN2 GA36_26(oper2[26], oper1[36], g36[26]);
AN2 GA36_27(oper2[27], oper1[36], g36[27]);
AN2 GA36_28(oper2[28], oper1[36], g36[28]);
AN2 GA36_29(oper2[29], oper1[36], g36[29]);
AN2 GA36_30(oper2[30], oper1[36], g36[30]);
AN2 GA36_31(oper2[31], oper1[36], g36[31]);
AN2 GA36_32(oper2[32], oper1[36], g36[32]);
AN2 GA36_33(oper2[33], oper1[36], g36[33]);
AN2 GA36_34(oper2[34], oper1[36], g36[34]);
AN2 GA36_35(oper2[35], oper1[36], g36[35]);
AN2 GA36_36(oper2[36], oper1[36], g36[36]);
AN2 GA36_37(oper2[37], oper1[36], g36[37]);
AN2 GA36_38(oper2[38], oper1[36], g36[38]);
AN2 GA36_39(oper2[39], oper1[36], g36[39]);
AN2 GA36_40(oper2[40], oper1[36], g36[40]);
AN2 GA36_41(oper2[41], oper1[36], g36[41]);
AN2 GA36_42(oper2[42], oper1[36], g36[42]);
AN2 GA36_43(oper2[43], oper1[36], g36[43]);
AN2 GA36_44(oper2[44], oper1[36], g36[44]);
AN2 GA36_45(oper2[45], oper1[36], g36[45]);
AN2 GA36_46(oper2[46], oper1[36], g36[46]);
AN2 GA36_47(oper2[47], oper1[36], g36[47]);
AN2 GA36_48(oper2[48], oper1[36], g36[48]);
AN2 GA36_49(oper2[49], oper1[36], g36[49]);
AN2 GA36_50(oper2[50], oper1[36], g36[50]);
AN2 GA36_51(oper2[51], oper1[36], g36[51]);
AN2 GA36_52(oper2[52], oper1[36], g36[52]);
AN2 GA36_53(oper2[53], oper1[36], g36[53]);
AN2 GA36_54(oper2[54], oper1[36], g36[54]);
AN2 GA36_55(oper2[55], oper1[36], g36[55]);
AN2 GA36_56(oper2[56], oper1[36], g36[56]);
AN2 GA36_57(oper2[57], oper1[36], g36[57]);
AN2 GA36_58(oper2[58], oper1[36], g36[58]);
AN2 GA36_59(oper2[59], oper1[36], g36[59]);
AN2 GA36_60(oper2[60], oper1[36], g36[60]);
AN2 GA36_61(oper2[61], oper1[36], g36[61]);
AN2 GA36_62(oper2[62], oper1[36], g36[62]);
AN2 GA36_63(oper2[63], oper1[36], g36[63]);
AN2 GA35_8(oper2[8], oper1[35], g35[8]);
AN2 GA35_9(oper2[9], oper1[35], g35[9]);
AN2 GA35_10(oper2[10], oper1[35], g35[10]);
AN2 GA35_11(oper2[11], oper1[35], g35[11]);
AN2 GA35_12(oper2[12], oper1[35], g35[12]);
AN2 GA35_13(oper2[13], oper1[35], g35[13]);
AN2 GA35_14(oper2[14], oper1[35], g35[14]);
AN2 GA35_15(oper2[15], oper1[35], g35[15]);
AN2 GA35_16(oper2[16], oper1[35], g35[16]);
AN2 GA35_17(oper2[17], oper1[35], g35[17]);
AN2 GA35_18(oper2[18], oper1[35], g35[18]);
AN2 GA35_19(oper2[19], oper1[35], g35[19]);
AN2 GA35_20(oper2[20], oper1[35], g35[20]);
AN2 GA35_21(oper2[21], oper1[35], g35[21]);
AN2 GA35_22(oper2[22], oper1[35], g35[22]);
AN2 GA35_23(oper2[23], oper1[35], g35[23]);
AN2 GA35_24(oper2[24], oper1[35], g35[24]);
AN2 GA35_25(oper2[25], oper1[35], g35[25]);
AN2 GA35_26(oper2[26], oper1[35], g35[26]);
AN2 GA35_27(oper2[27], oper1[35], g35[27]);
AN2 GA35_28(oper2[28], oper1[35], g35[28]);
AN2 GA35_29(oper2[29], oper1[35], g35[29]);
AN2 GA35_30(oper2[30], oper1[35], g35[30]);
AN2 GA35_31(oper2[31], oper1[35], g35[31]);
AN2 GA35_32(oper2[32], oper1[35], g35[32]);
AN2 GA35_33(oper2[33], oper1[35], g35[33]);
AN2 GA35_34(oper2[34], oper1[35], g35[34]);
AN2 GA35_35(oper2[35], oper1[35], g35[35]);
AN2 GA35_36(oper2[36], oper1[35], g35[36]);
AN2 GA35_37(oper2[37], oper1[35], g35[37]);
AN2 GA35_38(oper2[38], oper1[35], g35[38]);
AN2 GA35_39(oper2[39], oper1[35], g35[39]);
AN2 GA35_40(oper2[40], oper1[35], g35[40]);
AN2 GA35_41(oper2[41], oper1[35], g35[41]);
AN2 GA35_42(oper2[42], oper1[35], g35[42]);
AN2 GA35_43(oper2[43], oper1[35], g35[43]);
AN2 GA35_44(oper2[44], oper1[35], g35[44]);
AN2 GA35_45(oper2[45], oper1[35], g35[45]);
AN2 GA35_46(oper2[46], oper1[35], g35[46]);
AN2 GA35_47(oper2[47], oper1[35], g35[47]);
AN2 GA35_48(oper2[48], oper1[35], g35[48]);
AN2 GA35_49(oper2[49], oper1[35], g35[49]);
AN2 GA35_50(oper2[50], oper1[35], g35[50]);
AN2 GA35_51(oper2[51], oper1[35], g35[51]);
AN2 GA35_52(oper2[52], oper1[35], g35[52]);
AN2 GA35_53(oper2[53], oper1[35], g35[53]);
AN2 GA35_54(oper2[54], oper1[35], g35[54]);
AN2 GA35_55(oper2[55], oper1[35], g35[55]);
AN2 GA35_56(oper2[56], oper1[35], g35[56]);
AN2 GA35_57(oper2[57], oper1[35], g35[57]);
AN2 GA35_58(oper2[58], oper1[35], g35[58]);
AN2 GA35_59(oper2[59], oper1[35], g35[59]);
AN2 GA35_60(oper2[60], oper1[35], g35[60]);
AN2 GA35_61(oper2[61], oper1[35], g35[61]);
AN2 GA35_62(oper2[62], oper1[35], g35[62]);
AN2 GA35_63(oper2[63], oper1[35], g35[63]);
AN2 GA34_8(oper2[8], oper1[34], g34[8]);
AN2 GA34_9(oper2[9], oper1[34], g34[9]);
AN2 GA34_10(oper2[10], oper1[34], g34[10]);
AN2 GA34_11(oper2[11], oper1[34], g34[11]);
AN2 GA34_12(oper2[12], oper1[34], g34[12]);
AN2 GA34_13(oper2[13], oper1[34], g34[13]);
AN2 GA34_14(oper2[14], oper1[34], g34[14]);
AN2 GA34_15(oper2[15], oper1[34], g34[15]);
AN2 GA34_16(oper2[16], oper1[34], g34[16]);
AN2 GA34_17(oper2[17], oper1[34], g34[17]);
AN2 GA34_18(oper2[18], oper1[34], g34[18]);
AN2 GA34_19(oper2[19], oper1[34], g34[19]);
AN2 GA34_20(oper2[20], oper1[34], g34[20]);
AN2 GA34_21(oper2[21], oper1[34], g34[21]);
AN2 GA34_22(oper2[22], oper1[34], g34[22]);
AN2 GA34_23(oper2[23], oper1[34], g34[23]);
AN2 GA34_24(oper2[24], oper1[34], g34[24]);
AN2 GA34_25(oper2[25], oper1[34], g34[25]);
AN2 GA34_26(oper2[26], oper1[34], g34[26]);
AN2 GA34_27(oper2[27], oper1[34], g34[27]);
AN2 GA34_28(oper2[28], oper1[34], g34[28]);
AN2 GA34_29(oper2[29], oper1[34], g34[29]);
AN2 GA34_30(oper2[30], oper1[34], g34[30]);
AN2 GA34_31(oper2[31], oper1[34], g34[31]);
AN2 GA34_32(oper2[32], oper1[34], g34[32]);
AN2 GA34_33(oper2[33], oper1[34], g34[33]);
AN2 GA34_34(oper2[34], oper1[34], g34[34]);
AN2 GA34_35(oper2[35], oper1[34], g34[35]);
AN2 GA34_36(oper2[36], oper1[34], g34[36]);
AN2 GA34_37(oper2[37], oper1[34], g34[37]);
AN2 GA34_38(oper2[38], oper1[34], g34[38]);
AN2 GA34_39(oper2[39], oper1[34], g34[39]);
AN2 GA34_40(oper2[40], oper1[34], g34[40]);
AN2 GA34_41(oper2[41], oper1[34], g34[41]);
AN2 GA34_42(oper2[42], oper1[34], g34[42]);
AN2 GA34_43(oper2[43], oper1[34], g34[43]);
AN2 GA34_44(oper2[44], oper1[34], g34[44]);
AN2 GA34_45(oper2[45], oper1[34], g34[45]);
AN2 GA34_46(oper2[46], oper1[34], g34[46]);
AN2 GA34_47(oper2[47], oper1[34], g34[47]);
AN2 GA34_48(oper2[48], oper1[34], g34[48]);
AN2 GA34_49(oper2[49], oper1[34], g34[49]);
AN2 GA34_50(oper2[50], oper1[34], g34[50]);
AN2 GA34_51(oper2[51], oper1[34], g34[51]);
AN2 GA34_52(oper2[52], oper1[34], g34[52]);
AN2 GA34_53(oper2[53], oper1[34], g34[53]);
AN2 GA34_54(oper2[54], oper1[34], g34[54]);
AN2 GA34_55(oper2[55], oper1[34], g34[55]);
AN2 GA34_56(oper2[56], oper1[34], g34[56]);
AN2 GA34_57(oper2[57], oper1[34], g34[57]);
AN2 GA34_58(oper2[58], oper1[34], g34[58]);
AN2 GA34_59(oper2[59], oper1[34], g34[59]);
AN2 GA34_60(oper2[60], oper1[34], g34[60]);
AN2 GA34_61(oper2[61], oper1[34], g34[61]);
AN2 GA34_62(oper2[62], oper1[34], g34[62]);
AN2 GA34_63(oper2[63], oper1[34], g34[63]);
AN2 GA33_8(oper2[8], oper1[33], g33[8]);
AN2 GA33_9(oper2[9], oper1[33], g33[9]);
AN2 GA33_10(oper2[10], oper1[33], g33[10]);
AN2 GA33_11(oper2[11], oper1[33], g33[11]);
AN2 GA33_12(oper2[12], oper1[33], g33[12]);
AN2 GA33_13(oper2[13], oper1[33], g33[13]);
AN2 GA33_14(oper2[14], oper1[33], g33[14]);
AN2 GA33_15(oper2[15], oper1[33], g33[15]);
AN2 GA33_16(oper2[16], oper1[33], g33[16]);
AN2 GA33_17(oper2[17], oper1[33], g33[17]);
AN2 GA33_18(oper2[18], oper1[33], g33[18]);
AN2 GA33_19(oper2[19], oper1[33], g33[19]);
AN2 GA33_20(oper2[20], oper1[33], g33[20]);
AN2 GA33_21(oper2[21], oper1[33], g33[21]);
AN2 GA33_22(oper2[22], oper1[33], g33[22]);
AN2 GA33_23(oper2[23], oper1[33], g33[23]);
AN2 GA33_24(oper2[24], oper1[33], g33[24]);
AN2 GA33_25(oper2[25], oper1[33], g33[25]);
AN2 GA33_26(oper2[26], oper1[33], g33[26]);
AN2 GA33_27(oper2[27], oper1[33], g33[27]);
AN2 GA33_28(oper2[28], oper1[33], g33[28]);
AN2 GA33_29(oper2[29], oper1[33], g33[29]);
AN2 GA33_30(oper2[30], oper1[33], g33[30]);
AN2 GA33_31(oper2[31], oper1[33], g33[31]);
AN2 GA33_32(oper2[32], oper1[33], g33[32]);
AN2 GA33_33(oper2[33], oper1[33], g33[33]);
AN2 GA33_34(oper2[34], oper1[33], g33[34]);
AN2 GA33_35(oper2[35], oper1[33], g33[35]);
AN2 GA33_36(oper2[36], oper1[33], g33[36]);
AN2 GA33_37(oper2[37], oper1[33], g33[37]);
AN2 GA33_38(oper2[38], oper1[33], g33[38]);
AN2 GA33_39(oper2[39], oper1[33], g33[39]);
AN2 GA33_40(oper2[40], oper1[33], g33[40]);
AN2 GA33_41(oper2[41], oper1[33], g33[41]);
AN2 GA33_42(oper2[42], oper1[33], g33[42]);
AN2 GA33_43(oper2[43], oper1[33], g33[43]);
AN2 GA33_44(oper2[44], oper1[33], g33[44]);
AN2 GA33_45(oper2[45], oper1[33], g33[45]);
AN2 GA33_46(oper2[46], oper1[33], g33[46]);
AN2 GA33_47(oper2[47], oper1[33], g33[47]);
AN2 GA33_48(oper2[48], oper1[33], g33[48]);
AN2 GA33_49(oper2[49], oper1[33], g33[49]);
AN2 GA33_50(oper2[50], oper1[33], g33[50]);
AN2 GA33_51(oper2[51], oper1[33], g33[51]);
AN2 GA33_52(oper2[52], oper1[33], g33[52]);
AN2 GA33_53(oper2[53], oper1[33], g33[53]);
AN2 GA33_54(oper2[54], oper1[33], g33[54]);
AN2 GA33_55(oper2[55], oper1[33], g33[55]);
AN2 GA33_56(oper2[56], oper1[33], g33[56]);
AN2 GA33_57(oper2[57], oper1[33], g33[57]);
AN2 GA33_58(oper2[58], oper1[33], g33[58]);
AN2 GA33_59(oper2[59], oper1[33], g33[59]);
AN2 GA33_60(oper2[60], oper1[33], g33[60]);
AN2 GA33_61(oper2[61], oper1[33], g33[61]);
AN2 GA33_62(oper2[62], oper1[33], g33[62]);
AN2 GA33_63(oper2[63], oper1[33], g33[63]);
AN2 GA32_8(oper2[8], oper1[32], g32[8]);
AN2 GA32_9(oper2[9], oper1[32], g32[9]);
AN2 GA32_10(oper2[10], oper1[32], g32[10]);
AN2 GA32_11(oper2[11], oper1[32], g32[11]);
AN2 GA32_12(oper2[12], oper1[32], g32[12]);
AN2 GA32_13(oper2[13], oper1[32], g32[13]);
AN2 GA32_14(oper2[14], oper1[32], g32[14]);
AN2 GA32_15(oper2[15], oper1[32], g32[15]);
AN2 GA32_16(oper2[16], oper1[32], g32[16]);
AN2 GA32_17(oper2[17], oper1[32], g32[17]);
AN2 GA32_18(oper2[18], oper1[32], g32[18]);
AN2 GA32_19(oper2[19], oper1[32], g32[19]);
AN2 GA32_20(oper2[20], oper1[32], g32[20]);
AN2 GA32_21(oper2[21], oper1[32], g32[21]);
AN2 GA32_22(oper2[22], oper1[32], g32[22]);
AN2 GA32_23(oper2[23], oper1[32], g32[23]);
AN2 GA32_24(oper2[24], oper1[32], g32[24]);
AN2 GA32_25(oper2[25], oper1[32], g32[25]);
AN2 GA32_26(oper2[26], oper1[32], g32[26]);
AN2 GA32_27(oper2[27], oper1[32], g32[27]);
AN2 GA32_28(oper2[28], oper1[32], g32[28]);
AN2 GA32_29(oper2[29], oper1[32], g32[29]);
AN2 GA32_30(oper2[30], oper1[32], g32[30]);
AN2 GA32_31(oper2[31], oper1[32], g32[31]);
AN2 GA32_32(oper2[32], oper1[32], g32[32]);
AN2 GA32_33(oper2[33], oper1[32], g32[33]);
AN2 GA32_34(oper2[34], oper1[32], g32[34]);
AN2 GA32_35(oper2[35], oper1[32], g32[35]);
AN2 GA32_36(oper2[36], oper1[32], g32[36]);
AN2 GA32_37(oper2[37], oper1[32], g32[37]);
AN2 GA32_38(oper2[38], oper1[32], g32[38]);
AN2 GA32_39(oper2[39], oper1[32], g32[39]);
AN2 GA32_40(oper2[40], oper1[32], g32[40]);
AN2 GA32_41(oper2[41], oper1[32], g32[41]);
AN2 GA32_42(oper2[42], oper1[32], g32[42]);
AN2 GA32_43(oper2[43], oper1[32], g32[43]);
AN2 GA32_44(oper2[44], oper1[32], g32[44]);
AN2 GA32_45(oper2[45], oper1[32], g32[45]);
AN2 GA32_46(oper2[46], oper1[32], g32[46]);
AN2 GA32_47(oper2[47], oper1[32], g32[47]);
AN2 GA32_48(oper2[48], oper1[32], g32[48]);
AN2 GA32_49(oper2[49], oper1[32], g32[49]);
AN2 GA32_50(oper2[50], oper1[32], g32[50]);
AN2 GA32_51(oper2[51], oper1[32], g32[51]);
AN2 GA32_52(oper2[52], oper1[32], g32[52]);
AN2 GA32_53(oper2[53], oper1[32], g32[53]);
AN2 GA32_54(oper2[54], oper1[32], g32[54]);
AN2 GA32_55(oper2[55], oper1[32], g32[55]);
AN2 GA32_56(oper2[56], oper1[32], g32[56]);
AN2 GA32_57(oper2[57], oper1[32], g32[57]);
AN2 GA32_58(oper2[58], oper1[32], g32[58]);
AN2 GA32_59(oper2[59], oper1[32], g32[59]);
AN2 GA32_60(oper2[60], oper1[32], g32[60]);
AN2 GA32_61(oper2[61], oper1[32], g32[61]);
AN2 GA32_62(oper2[62], oper1[32], g32[62]);
AN2 GA32_63(oper2[63], oper1[32], g32[63]);
AN2 GA31_8(oper2[8], oper1[31], g31[8]);
AN2 GA31_9(oper2[9], oper1[31], g31[9]);
AN2 GA31_10(oper2[10], oper1[31], g31[10]);
AN2 GA31_11(oper2[11], oper1[31], g31[11]);
AN2 GA31_12(oper2[12], oper1[31], g31[12]);
AN2 GA31_13(oper2[13], oper1[31], g31[13]);
AN2 GA31_14(oper2[14], oper1[31], g31[14]);
AN2 GA31_15(oper2[15], oper1[31], g31[15]);
AN2 GA31_16(oper2[16], oper1[31], g31[16]);
AN2 GA31_17(oper2[17], oper1[31], g31[17]);
AN2 GA31_18(oper2[18], oper1[31], g31[18]);
AN2 GA31_19(oper2[19], oper1[31], g31[19]);
AN2 GA31_20(oper2[20], oper1[31], g31[20]);
AN2 GA31_21(oper2[21], oper1[31], g31[21]);
AN2 GA31_22(oper2[22], oper1[31], g31[22]);
AN2 GA31_23(oper2[23], oper1[31], g31[23]);
AN2 GA31_24(oper2[24], oper1[31], g31[24]);
AN2 GA31_25(oper2[25], oper1[31], g31[25]);
AN2 GA31_26(oper2[26], oper1[31], g31[26]);
AN2 GA31_27(oper2[27], oper1[31], g31[27]);
AN2 GA31_28(oper2[28], oper1[31], g31[28]);
AN2 GA31_29(oper2[29], oper1[31], g31[29]);
AN2 GA31_30(oper2[30], oper1[31], g31[30]);
AN2 GA31_31(oper2[31], oper1[31], g31[31]);
AN2 GA31_32(oper2[32], oper1[31], g31[32]);
AN2 GA31_33(oper2[33], oper1[31], g31[33]);
AN2 GA31_34(oper2[34], oper1[31], g31[34]);
AN2 GA31_35(oper2[35], oper1[31], g31[35]);
AN2 GA31_36(oper2[36], oper1[31], g31[36]);
AN2 GA31_37(oper2[37], oper1[31], g31[37]);
AN2 GA31_38(oper2[38], oper1[31], g31[38]);
AN2 GA31_39(oper2[39], oper1[31], g31[39]);
AN2 GA31_40(oper2[40], oper1[31], g31[40]);
AN2 GA31_41(oper2[41], oper1[31], g31[41]);
AN2 GA31_42(oper2[42], oper1[31], g31[42]);
AN2 GA31_43(oper2[43], oper1[31], g31[43]);
AN2 GA31_44(oper2[44], oper1[31], g31[44]);
AN2 GA31_45(oper2[45], oper1[31], g31[45]);
AN2 GA31_46(oper2[46], oper1[31], g31[46]);
AN2 GA31_47(oper2[47], oper1[31], g31[47]);
AN2 GA31_48(oper2[48], oper1[31], g31[48]);
AN2 GA31_49(oper2[49], oper1[31], g31[49]);
AN2 GA31_50(oper2[50], oper1[31], g31[50]);
AN2 GA31_51(oper2[51], oper1[31], g31[51]);
AN2 GA31_52(oper2[52], oper1[31], g31[52]);
AN2 GA31_53(oper2[53], oper1[31], g31[53]);
AN2 GA31_54(oper2[54], oper1[31], g31[54]);
AN2 GA31_55(oper2[55], oper1[31], g31[55]);
AN2 GA31_56(oper2[56], oper1[31], g31[56]);
AN2 GA31_57(oper2[57], oper1[31], g31[57]);
AN2 GA31_58(oper2[58], oper1[31], g31[58]);
AN2 GA31_59(oper2[59], oper1[31], g31[59]);
AN2 GA31_60(oper2[60], oper1[31], g31[60]);
AN2 GA31_61(oper2[61], oper1[31], g31[61]);
AN2 GA31_62(oper2[62], oper1[31], g31[62]);
AN2 GA31_63(oper2[63], oper1[31], g31[63]);
AN2 GA30_8(oper2[8], oper1[30], g30[8]);
AN2 GA30_9(oper2[9], oper1[30], g30[9]);
AN2 GA30_10(oper2[10], oper1[30], g30[10]);
AN2 GA30_11(oper2[11], oper1[30], g30[11]);
AN2 GA30_12(oper2[12], oper1[30], g30[12]);
AN2 GA30_13(oper2[13], oper1[30], g30[13]);
AN2 GA30_14(oper2[14], oper1[30], g30[14]);
AN2 GA30_15(oper2[15], oper1[30], g30[15]);
AN2 GA30_16(oper2[16], oper1[30], g30[16]);
AN2 GA30_17(oper2[17], oper1[30], g30[17]);
AN2 GA30_18(oper2[18], oper1[30], g30[18]);
AN2 GA30_19(oper2[19], oper1[30], g30[19]);
AN2 GA30_20(oper2[20], oper1[30], g30[20]);
AN2 GA30_21(oper2[21], oper1[30], g30[21]);
AN2 GA30_22(oper2[22], oper1[30], g30[22]);
AN2 GA30_23(oper2[23], oper1[30], g30[23]);
AN2 GA30_24(oper2[24], oper1[30], g30[24]);
AN2 GA30_25(oper2[25], oper1[30], g30[25]);
AN2 GA30_26(oper2[26], oper1[30], g30[26]);
AN2 GA30_27(oper2[27], oper1[30], g30[27]);
AN2 GA30_28(oper2[28], oper1[30], g30[28]);
AN2 GA30_29(oper2[29], oper1[30], g30[29]);
AN2 GA30_30(oper2[30], oper1[30], g30[30]);
AN2 GA30_31(oper2[31], oper1[30], g30[31]);
AN2 GA30_32(oper2[32], oper1[30], g30[32]);
AN2 GA30_33(oper2[33], oper1[30], g30[33]);
AN2 GA30_34(oper2[34], oper1[30], g30[34]);
AN2 GA30_35(oper2[35], oper1[30], g30[35]);
AN2 GA30_36(oper2[36], oper1[30], g30[36]);
AN2 GA30_37(oper2[37], oper1[30], g30[37]);
AN2 GA30_38(oper2[38], oper1[30], g30[38]);
AN2 GA30_39(oper2[39], oper1[30], g30[39]);
AN2 GA30_40(oper2[40], oper1[30], g30[40]);
AN2 GA30_41(oper2[41], oper1[30], g30[41]);
AN2 GA30_42(oper2[42], oper1[30], g30[42]);
AN2 GA30_43(oper2[43], oper1[30], g30[43]);
AN2 GA30_44(oper2[44], oper1[30], g30[44]);
AN2 GA30_45(oper2[45], oper1[30], g30[45]);
AN2 GA30_46(oper2[46], oper1[30], g30[46]);
AN2 GA30_47(oper2[47], oper1[30], g30[47]);
AN2 GA30_48(oper2[48], oper1[30], g30[48]);
AN2 GA30_49(oper2[49], oper1[30], g30[49]);
AN2 GA30_50(oper2[50], oper1[30], g30[50]);
AN2 GA30_51(oper2[51], oper1[30], g30[51]);
AN2 GA30_52(oper2[52], oper1[30], g30[52]);
AN2 GA30_53(oper2[53], oper1[30], g30[53]);
AN2 GA30_54(oper2[54], oper1[30], g30[54]);
AN2 GA30_55(oper2[55], oper1[30], g30[55]);
AN2 GA30_56(oper2[56], oper1[30], g30[56]);
AN2 GA30_57(oper2[57], oper1[30], g30[57]);
AN2 GA30_58(oper2[58], oper1[30], g30[58]);
AN2 GA30_59(oper2[59], oper1[30], g30[59]);
AN2 GA30_60(oper2[60], oper1[30], g30[60]);
AN2 GA30_61(oper2[61], oper1[30], g30[61]);
AN2 GA30_62(oper2[62], oper1[30], g30[62]);
AN2 GA30_63(oper2[63], oper1[30], g30[63]);
AN2 GA29_8(oper2[8], oper1[29], g29[8]);
AN2 GA29_9(oper2[9], oper1[29], g29[9]);
AN2 GA29_10(oper2[10], oper1[29], g29[10]);
AN2 GA29_11(oper2[11], oper1[29], g29[11]);
AN2 GA29_12(oper2[12], oper1[29], g29[12]);
AN2 GA29_13(oper2[13], oper1[29], g29[13]);
AN2 GA29_14(oper2[14], oper1[29], g29[14]);
AN2 GA29_15(oper2[15], oper1[29], g29[15]);
AN2 GA29_16(oper2[16], oper1[29], g29[16]);
AN2 GA29_17(oper2[17], oper1[29], g29[17]);
AN2 GA29_18(oper2[18], oper1[29], g29[18]);
AN2 GA29_19(oper2[19], oper1[29], g29[19]);
AN2 GA29_20(oper2[20], oper1[29], g29[20]);
AN2 GA29_21(oper2[21], oper1[29], g29[21]);
AN2 GA29_22(oper2[22], oper1[29], g29[22]);
AN2 GA29_23(oper2[23], oper1[29], g29[23]);
AN2 GA29_24(oper2[24], oper1[29], g29[24]);
AN2 GA29_25(oper2[25], oper1[29], g29[25]);
AN2 GA29_26(oper2[26], oper1[29], g29[26]);
AN2 GA29_27(oper2[27], oper1[29], g29[27]);
AN2 GA29_28(oper2[28], oper1[29], g29[28]);
AN2 GA29_29(oper2[29], oper1[29], g29[29]);
AN2 GA29_30(oper2[30], oper1[29], g29[30]);
AN2 GA29_31(oper2[31], oper1[29], g29[31]);
AN2 GA29_32(oper2[32], oper1[29], g29[32]);
AN2 GA29_33(oper2[33], oper1[29], g29[33]);
AN2 GA29_34(oper2[34], oper1[29], g29[34]);
AN2 GA29_35(oper2[35], oper1[29], g29[35]);
AN2 GA29_36(oper2[36], oper1[29], g29[36]);
AN2 GA29_37(oper2[37], oper1[29], g29[37]);
AN2 GA29_38(oper2[38], oper1[29], g29[38]);
AN2 GA29_39(oper2[39], oper1[29], g29[39]);
AN2 GA29_40(oper2[40], oper1[29], g29[40]);
AN2 GA29_41(oper2[41], oper1[29], g29[41]);
AN2 GA29_42(oper2[42], oper1[29], g29[42]);
AN2 GA29_43(oper2[43], oper1[29], g29[43]);
AN2 GA29_44(oper2[44], oper1[29], g29[44]);
AN2 GA29_45(oper2[45], oper1[29], g29[45]);
AN2 GA29_46(oper2[46], oper1[29], g29[46]);
AN2 GA29_47(oper2[47], oper1[29], g29[47]);
AN2 GA29_48(oper2[48], oper1[29], g29[48]);
AN2 GA29_49(oper2[49], oper1[29], g29[49]);
AN2 GA29_50(oper2[50], oper1[29], g29[50]);
AN2 GA29_51(oper2[51], oper1[29], g29[51]);
AN2 GA29_52(oper2[52], oper1[29], g29[52]);
AN2 GA29_53(oper2[53], oper1[29], g29[53]);
AN2 GA29_54(oper2[54], oper1[29], g29[54]);
AN2 GA29_55(oper2[55], oper1[29], g29[55]);
AN2 GA29_56(oper2[56], oper1[29], g29[56]);
AN2 GA29_57(oper2[57], oper1[29], g29[57]);
AN2 GA29_58(oper2[58], oper1[29], g29[58]);
AN2 GA29_59(oper2[59], oper1[29], g29[59]);
AN2 GA29_60(oper2[60], oper1[29], g29[60]);
AN2 GA29_61(oper2[61], oper1[29], g29[61]);
AN2 GA29_62(oper2[62], oper1[29], g29[62]);
AN2 GA29_63(oper2[63], oper1[29], g29[63]);
AN2 GA28_8(oper2[8], oper1[28], g28[8]);
AN2 GA28_9(oper2[9], oper1[28], g28[9]);
AN2 GA28_10(oper2[10], oper1[28], g28[10]);
AN2 GA28_11(oper2[11], oper1[28], g28[11]);
AN2 GA28_12(oper2[12], oper1[28], g28[12]);
AN2 GA28_13(oper2[13], oper1[28], g28[13]);
AN2 GA28_14(oper2[14], oper1[28], g28[14]);
AN2 GA28_15(oper2[15], oper1[28], g28[15]);
AN2 GA28_16(oper2[16], oper1[28], g28[16]);
AN2 GA28_17(oper2[17], oper1[28], g28[17]);
AN2 GA28_18(oper2[18], oper1[28], g28[18]);
AN2 GA28_19(oper2[19], oper1[28], g28[19]);
AN2 GA28_20(oper2[20], oper1[28], g28[20]);
AN2 GA28_21(oper2[21], oper1[28], g28[21]);
AN2 GA28_22(oper2[22], oper1[28], g28[22]);
AN2 GA28_23(oper2[23], oper1[28], g28[23]);
AN2 GA28_24(oper2[24], oper1[28], g28[24]);
AN2 GA28_25(oper2[25], oper1[28], g28[25]);
AN2 GA28_26(oper2[26], oper1[28], g28[26]);
AN2 GA28_27(oper2[27], oper1[28], g28[27]);
AN2 GA28_28(oper2[28], oper1[28], g28[28]);
AN2 GA28_29(oper2[29], oper1[28], g28[29]);
AN2 GA28_30(oper2[30], oper1[28], g28[30]);
AN2 GA28_31(oper2[31], oper1[28], g28[31]);
AN2 GA28_32(oper2[32], oper1[28], g28[32]);
AN2 GA28_33(oper2[33], oper1[28], g28[33]);
AN2 GA28_34(oper2[34], oper1[28], g28[34]);
AN2 GA28_35(oper2[35], oper1[28], g28[35]);
AN2 GA28_36(oper2[36], oper1[28], g28[36]);
AN2 GA28_37(oper2[37], oper1[28], g28[37]);
AN2 GA28_38(oper2[38], oper1[28], g28[38]);
AN2 GA28_39(oper2[39], oper1[28], g28[39]);
AN2 GA28_40(oper2[40], oper1[28], g28[40]);
AN2 GA28_41(oper2[41], oper1[28], g28[41]);
AN2 GA28_42(oper2[42], oper1[28], g28[42]);
AN2 GA28_43(oper2[43], oper1[28], g28[43]);
AN2 GA28_44(oper2[44], oper1[28], g28[44]);
AN2 GA28_45(oper2[45], oper1[28], g28[45]);
AN2 GA28_46(oper2[46], oper1[28], g28[46]);
AN2 GA28_47(oper2[47], oper1[28], g28[47]);
AN2 GA28_48(oper2[48], oper1[28], g28[48]);
AN2 GA28_49(oper2[49], oper1[28], g28[49]);
AN2 GA28_50(oper2[50], oper1[28], g28[50]);
AN2 GA28_51(oper2[51], oper1[28], g28[51]);
AN2 GA28_52(oper2[52], oper1[28], g28[52]);
AN2 GA28_53(oper2[53], oper1[28], g28[53]);
AN2 GA28_54(oper2[54], oper1[28], g28[54]);
AN2 GA28_55(oper2[55], oper1[28], g28[55]);
AN2 GA28_56(oper2[56], oper1[28], g28[56]);
AN2 GA28_57(oper2[57], oper1[28], g28[57]);
AN2 GA28_58(oper2[58], oper1[28], g28[58]);
AN2 GA28_59(oper2[59], oper1[28], g28[59]);
AN2 GA28_60(oper2[60], oper1[28], g28[60]);
AN2 GA28_61(oper2[61], oper1[28], g28[61]);
AN2 GA28_62(oper2[62], oper1[28], g28[62]);
AN2 GA28_63(oper2[63], oper1[28], g28[63]);
AN2 GA27_8(oper2[8], oper1[27], g27[8]);
AN2 GA27_9(oper2[9], oper1[27], g27[9]);
AN2 GA27_10(oper2[10], oper1[27], g27[10]);
AN2 GA27_11(oper2[11], oper1[27], g27[11]);
AN2 GA27_12(oper2[12], oper1[27], g27[12]);
AN2 GA27_13(oper2[13], oper1[27], g27[13]);
AN2 GA27_14(oper2[14], oper1[27], g27[14]);
AN2 GA27_15(oper2[15], oper1[27], g27[15]);
AN2 GA27_16(oper2[16], oper1[27], g27[16]);
AN2 GA27_17(oper2[17], oper1[27], g27[17]);
AN2 GA27_18(oper2[18], oper1[27], g27[18]);
AN2 GA27_19(oper2[19], oper1[27], g27[19]);
AN2 GA27_20(oper2[20], oper1[27], g27[20]);
AN2 GA27_21(oper2[21], oper1[27], g27[21]);
AN2 GA27_22(oper2[22], oper1[27], g27[22]);
AN2 GA27_23(oper2[23], oper1[27], g27[23]);
AN2 GA27_24(oper2[24], oper1[27], g27[24]);
AN2 GA27_25(oper2[25], oper1[27], g27[25]);
AN2 GA27_26(oper2[26], oper1[27], g27[26]);
AN2 GA27_27(oper2[27], oper1[27], g27[27]);
AN2 GA27_28(oper2[28], oper1[27], g27[28]);
AN2 GA27_29(oper2[29], oper1[27], g27[29]);
AN2 GA27_30(oper2[30], oper1[27], g27[30]);
AN2 GA27_31(oper2[31], oper1[27], g27[31]);
AN2 GA27_32(oper2[32], oper1[27], g27[32]);
AN2 GA27_33(oper2[33], oper1[27], g27[33]);
AN2 GA27_34(oper2[34], oper1[27], g27[34]);
AN2 GA27_35(oper2[35], oper1[27], g27[35]);
AN2 GA27_36(oper2[36], oper1[27], g27[36]);
AN2 GA27_37(oper2[37], oper1[27], g27[37]);
AN2 GA27_38(oper2[38], oper1[27], g27[38]);
AN2 GA27_39(oper2[39], oper1[27], g27[39]);
AN2 GA27_40(oper2[40], oper1[27], g27[40]);
AN2 GA27_41(oper2[41], oper1[27], g27[41]);
AN2 GA27_42(oper2[42], oper1[27], g27[42]);
AN2 GA27_43(oper2[43], oper1[27], g27[43]);
AN2 GA27_44(oper2[44], oper1[27], g27[44]);
AN2 GA27_45(oper2[45], oper1[27], g27[45]);
AN2 GA27_46(oper2[46], oper1[27], g27[46]);
AN2 GA27_47(oper2[47], oper1[27], g27[47]);
AN2 GA27_48(oper2[48], oper1[27], g27[48]);
AN2 GA27_49(oper2[49], oper1[27], g27[49]);
AN2 GA27_50(oper2[50], oper1[27], g27[50]);
AN2 GA27_51(oper2[51], oper1[27], g27[51]);
AN2 GA27_52(oper2[52], oper1[27], g27[52]);
AN2 GA27_53(oper2[53], oper1[27], g27[53]);
AN2 GA27_54(oper2[54], oper1[27], g27[54]);
AN2 GA27_55(oper2[55], oper1[27], g27[55]);
AN2 GA27_56(oper2[56], oper1[27], g27[56]);
AN2 GA27_57(oper2[57], oper1[27], g27[57]);
AN2 GA27_58(oper2[58], oper1[27], g27[58]);
AN2 GA27_59(oper2[59], oper1[27], g27[59]);
AN2 GA27_60(oper2[60], oper1[27], g27[60]);
AN2 GA27_61(oper2[61], oper1[27], g27[61]);
AN2 GA27_62(oper2[62], oper1[27], g27[62]);
AN2 GA27_63(oper2[63], oper1[27], g27[63]);
AN2 GA26_8(oper2[8], oper1[26], g26[8]);
AN2 GA26_9(oper2[9], oper1[26], g26[9]);
AN2 GA26_10(oper2[10], oper1[26], g26[10]);
AN2 GA26_11(oper2[11], oper1[26], g26[11]);
AN2 GA26_12(oper2[12], oper1[26], g26[12]);
AN2 GA26_13(oper2[13], oper1[26], g26[13]);
AN2 GA26_14(oper2[14], oper1[26], g26[14]);
AN2 GA26_15(oper2[15], oper1[26], g26[15]);
AN2 GA26_16(oper2[16], oper1[26], g26[16]);
AN2 GA26_17(oper2[17], oper1[26], g26[17]);
AN2 GA26_18(oper2[18], oper1[26], g26[18]);
AN2 GA26_19(oper2[19], oper1[26], g26[19]);
AN2 GA26_20(oper2[20], oper1[26], g26[20]);
AN2 GA26_21(oper2[21], oper1[26], g26[21]);
AN2 GA26_22(oper2[22], oper1[26], g26[22]);
AN2 GA26_23(oper2[23], oper1[26], g26[23]);
AN2 GA26_24(oper2[24], oper1[26], g26[24]);
AN2 GA26_25(oper2[25], oper1[26], g26[25]);
AN2 GA26_26(oper2[26], oper1[26], g26[26]);
AN2 GA26_27(oper2[27], oper1[26], g26[27]);
AN2 GA26_28(oper2[28], oper1[26], g26[28]);
AN2 GA26_29(oper2[29], oper1[26], g26[29]);
AN2 GA26_30(oper2[30], oper1[26], g26[30]);
AN2 GA26_31(oper2[31], oper1[26], g26[31]);
AN2 GA26_32(oper2[32], oper1[26], g26[32]);
AN2 GA26_33(oper2[33], oper1[26], g26[33]);
AN2 GA26_34(oper2[34], oper1[26], g26[34]);
AN2 GA26_35(oper2[35], oper1[26], g26[35]);
AN2 GA26_36(oper2[36], oper1[26], g26[36]);
AN2 GA26_37(oper2[37], oper1[26], g26[37]);
AN2 GA26_38(oper2[38], oper1[26], g26[38]);
AN2 GA26_39(oper2[39], oper1[26], g26[39]);
AN2 GA26_40(oper2[40], oper1[26], g26[40]);
AN2 GA26_41(oper2[41], oper1[26], g26[41]);
AN2 GA26_42(oper2[42], oper1[26], g26[42]);
AN2 GA26_43(oper2[43], oper1[26], g26[43]);
AN2 GA26_44(oper2[44], oper1[26], g26[44]);
AN2 GA26_45(oper2[45], oper1[26], g26[45]);
AN2 GA26_46(oper2[46], oper1[26], g26[46]);
AN2 GA26_47(oper2[47], oper1[26], g26[47]);
AN2 GA26_48(oper2[48], oper1[26], g26[48]);
AN2 GA26_49(oper2[49], oper1[26], g26[49]);
AN2 GA26_50(oper2[50], oper1[26], g26[50]);
AN2 GA26_51(oper2[51], oper1[26], g26[51]);
AN2 GA26_52(oper2[52], oper1[26], g26[52]);
AN2 GA26_53(oper2[53], oper1[26], g26[53]);
AN2 GA26_54(oper2[54], oper1[26], g26[54]);
AN2 GA26_55(oper2[55], oper1[26], g26[55]);
AN2 GA26_56(oper2[56], oper1[26], g26[56]);
AN2 GA26_57(oper2[57], oper1[26], g26[57]);
AN2 GA26_58(oper2[58], oper1[26], g26[58]);
AN2 GA26_59(oper2[59], oper1[26], g26[59]);
AN2 GA26_60(oper2[60], oper1[26], g26[60]);
AN2 GA26_61(oper2[61], oper1[26], g26[61]);
AN2 GA26_62(oper2[62], oper1[26], g26[62]);
AN2 GA26_63(oper2[63], oper1[26], g26[63]);
AN2 GA25_8(oper2[8], oper1[25], g25[8]);
AN2 GA25_9(oper2[9], oper1[25], g25[9]);
AN2 GA25_10(oper2[10], oper1[25], g25[10]);
AN2 GA25_11(oper2[11], oper1[25], g25[11]);
AN2 GA25_12(oper2[12], oper1[25], g25[12]);
AN2 GA25_13(oper2[13], oper1[25], g25[13]);
AN2 GA25_14(oper2[14], oper1[25], g25[14]);
AN2 GA25_15(oper2[15], oper1[25], g25[15]);
AN2 GA25_16(oper2[16], oper1[25], g25[16]);
AN2 GA25_17(oper2[17], oper1[25], g25[17]);
AN2 GA25_18(oper2[18], oper1[25], g25[18]);
AN2 GA25_19(oper2[19], oper1[25], g25[19]);
AN2 GA25_20(oper2[20], oper1[25], g25[20]);
AN2 GA25_21(oper2[21], oper1[25], g25[21]);
AN2 GA25_22(oper2[22], oper1[25], g25[22]);
AN2 GA25_23(oper2[23], oper1[25], g25[23]);
AN2 GA25_24(oper2[24], oper1[25], g25[24]);
AN2 GA25_25(oper2[25], oper1[25], g25[25]);
AN2 GA25_26(oper2[26], oper1[25], g25[26]);
AN2 GA25_27(oper2[27], oper1[25], g25[27]);
AN2 GA25_28(oper2[28], oper1[25], g25[28]);
AN2 GA25_29(oper2[29], oper1[25], g25[29]);
AN2 GA25_30(oper2[30], oper1[25], g25[30]);
AN2 GA25_31(oper2[31], oper1[25], g25[31]);
AN2 GA25_32(oper2[32], oper1[25], g25[32]);
AN2 GA25_33(oper2[33], oper1[25], g25[33]);
AN2 GA25_34(oper2[34], oper1[25], g25[34]);
AN2 GA25_35(oper2[35], oper1[25], g25[35]);
AN2 GA25_36(oper2[36], oper1[25], g25[36]);
AN2 GA25_37(oper2[37], oper1[25], g25[37]);
AN2 GA25_38(oper2[38], oper1[25], g25[38]);
AN2 GA25_39(oper2[39], oper1[25], g25[39]);
AN2 GA25_40(oper2[40], oper1[25], g25[40]);
AN2 GA25_41(oper2[41], oper1[25], g25[41]);
AN2 GA25_42(oper2[42], oper1[25], g25[42]);
AN2 GA25_43(oper2[43], oper1[25], g25[43]);
AN2 GA25_44(oper2[44], oper1[25], g25[44]);
AN2 GA25_45(oper2[45], oper1[25], g25[45]);
AN2 GA25_46(oper2[46], oper1[25], g25[46]);
AN2 GA25_47(oper2[47], oper1[25], g25[47]);
AN2 GA25_48(oper2[48], oper1[25], g25[48]);
AN2 GA25_49(oper2[49], oper1[25], g25[49]);
AN2 GA25_50(oper2[50], oper1[25], g25[50]);
AN2 GA25_51(oper2[51], oper1[25], g25[51]);
AN2 GA25_52(oper2[52], oper1[25], g25[52]);
AN2 GA25_53(oper2[53], oper1[25], g25[53]);
AN2 GA25_54(oper2[54], oper1[25], g25[54]);
AN2 GA25_55(oper2[55], oper1[25], g25[55]);
AN2 GA25_56(oper2[56], oper1[25], g25[56]);
AN2 GA25_57(oper2[57], oper1[25], g25[57]);
AN2 GA25_58(oper2[58], oper1[25], g25[58]);
AN2 GA25_59(oper2[59], oper1[25], g25[59]);
AN2 GA25_60(oper2[60], oper1[25], g25[60]);
AN2 GA25_61(oper2[61], oper1[25], g25[61]);
AN2 GA25_62(oper2[62], oper1[25], g25[62]);
AN2 GA25_63(oper2[63], oper1[25], g25[63]);
AN2 GA24_8(oper2[8], oper1[24], g24[8]);
AN2 GA24_9(oper2[9], oper1[24], g24[9]);
AN2 GA24_10(oper2[10], oper1[24], g24[10]);
AN2 GA24_11(oper2[11], oper1[24], g24[11]);
AN2 GA24_12(oper2[12], oper1[24], g24[12]);
AN2 GA24_13(oper2[13], oper1[24], g24[13]);
AN2 GA24_14(oper2[14], oper1[24], g24[14]);
AN2 GA24_15(oper2[15], oper1[24], g24[15]);
AN2 GA24_16(oper2[16], oper1[24], g24[16]);
AN2 GA24_17(oper2[17], oper1[24], g24[17]);
AN2 GA24_18(oper2[18], oper1[24], g24[18]);
AN2 GA24_19(oper2[19], oper1[24], g24[19]);
AN2 GA24_20(oper2[20], oper1[24], g24[20]);
AN2 GA24_21(oper2[21], oper1[24], g24[21]);
AN2 GA24_22(oper2[22], oper1[24], g24[22]);
AN2 GA24_23(oper2[23], oper1[24], g24[23]);
AN2 GA24_24(oper2[24], oper1[24], g24[24]);
AN2 GA24_25(oper2[25], oper1[24], g24[25]);
AN2 GA24_26(oper2[26], oper1[24], g24[26]);
AN2 GA24_27(oper2[27], oper1[24], g24[27]);
AN2 GA24_28(oper2[28], oper1[24], g24[28]);
AN2 GA24_29(oper2[29], oper1[24], g24[29]);
AN2 GA24_30(oper2[30], oper1[24], g24[30]);
AN2 GA24_31(oper2[31], oper1[24], g24[31]);
AN2 GA24_32(oper2[32], oper1[24], g24[32]);
AN2 GA24_33(oper2[33], oper1[24], g24[33]);
AN2 GA24_34(oper2[34], oper1[24], g24[34]);
AN2 GA24_35(oper2[35], oper1[24], g24[35]);
AN2 GA24_36(oper2[36], oper1[24], g24[36]);
AN2 GA24_37(oper2[37], oper1[24], g24[37]);
AN2 GA24_38(oper2[38], oper1[24], g24[38]);
AN2 GA24_39(oper2[39], oper1[24], g24[39]);
AN2 GA24_40(oper2[40], oper1[24], g24[40]);
AN2 GA24_41(oper2[41], oper1[24], g24[41]);
AN2 GA24_42(oper2[42], oper1[24], g24[42]);
AN2 GA24_43(oper2[43], oper1[24], g24[43]);
AN2 GA24_44(oper2[44], oper1[24], g24[44]);
AN2 GA24_45(oper2[45], oper1[24], g24[45]);
AN2 GA24_46(oper2[46], oper1[24], g24[46]);
AN2 GA24_47(oper2[47], oper1[24], g24[47]);
AN2 GA24_48(oper2[48], oper1[24], g24[48]);
AN2 GA24_49(oper2[49], oper1[24], g24[49]);
AN2 GA24_50(oper2[50], oper1[24], g24[50]);
AN2 GA24_51(oper2[51], oper1[24], g24[51]);
AN2 GA24_52(oper2[52], oper1[24], g24[52]);
AN2 GA24_53(oper2[53], oper1[24], g24[53]);
AN2 GA24_54(oper2[54], oper1[24], g24[54]);
AN2 GA24_55(oper2[55], oper1[24], g24[55]);
AN2 GA24_56(oper2[56], oper1[24], g24[56]);
AN2 GA24_57(oper2[57], oper1[24], g24[57]);
AN2 GA24_58(oper2[58], oper1[24], g24[58]);
AN2 GA24_59(oper2[59], oper1[24], g24[59]);
AN2 GA24_60(oper2[60], oper1[24], g24[60]);
AN2 GA24_61(oper2[61], oper1[24], g24[61]);
AN2 GA24_62(oper2[62], oper1[24], g24[62]);
AN2 GA24_63(oper2[63], oper1[24], g24[63]);
AN2 GA23_8(oper2[8], oper1[23], g23[8]);
AN2 GA23_9(oper2[9], oper1[23], g23[9]);
AN2 GA23_10(oper2[10], oper1[23], g23[10]);
AN2 GA23_11(oper2[11], oper1[23], g23[11]);
AN2 GA23_12(oper2[12], oper1[23], g23[12]);
AN2 GA23_13(oper2[13], oper1[23], g23[13]);
AN2 GA23_14(oper2[14], oper1[23], g23[14]);
AN2 GA23_15(oper2[15], oper1[23], g23[15]);
AN2 GA23_16(oper2[16], oper1[23], g23[16]);
AN2 GA23_17(oper2[17], oper1[23], g23[17]);
AN2 GA23_18(oper2[18], oper1[23], g23[18]);
AN2 GA23_19(oper2[19], oper1[23], g23[19]);
AN2 GA23_20(oper2[20], oper1[23], g23[20]);
AN2 GA23_21(oper2[21], oper1[23], g23[21]);
AN2 GA23_22(oper2[22], oper1[23], g23[22]);
AN2 GA23_23(oper2[23], oper1[23], g23[23]);
AN2 GA23_24(oper2[24], oper1[23], g23[24]);
AN2 GA23_25(oper2[25], oper1[23], g23[25]);
AN2 GA23_26(oper2[26], oper1[23], g23[26]);
AN2 GA23_27(oper2[27], oper1[23], g23[27]);
AN2 GA23_28(oper2[28], oper1[23], g23[28]);
AN2 GA23_29(oper2[29], oper1[23], g23[29]);
AN2 GA23_30(oper2[30], oper1[23], g23[30]);
AN2 GA23_31(oper2[31], oper1[23], g23[31]);
AN2 GA23_32(oper2[32], oper1[23], g23[32]);
AN2 GA23_33(oper2[33], oper1[23], g23[33]);
AN2 GA23_34(oper2[34], oper1[23], g23[34]);
AN2 GA23_35(oper2[35], oper1[23], g23[35]);
AN2 GA23_36(oper2[36], oper1[23], g23[36]);
AN2 GA23_37(oper2[37], oper1[23], g23[37]);
AN2 GA23_38(oper2[38], oper1[23], g23[38]);
AN2 GA23_39(oper2[39], oper1[23], g23[39]);
AN2 GA23_40(oper2[40], oper1[23], g23[40]);
AN2 GA23_41(oper2[41], oper1[23], g23[41]);
AN2 GA23_42(oper2[42], oper1[23], g23[42]);
AN2 GA23_43(oper2[43], oper1[23], g23[43]);
AN2 GA23_44(oper2[44], oper1[23], g23[44]);
AN2 GA23_45(oper2[45], oper1[23], g23[45]);
AN2 GA23_46(oper2[46], oper1[23], g23[46]);
AN2 GA23_47(oper2[47], oper1[23], g23[47]);
AN2 GA23_48(oper2[48], oper1[23], g23[48]);
AN2 GA23_49(oper2[49], oper1[23], g23[49]);
AN2 GA23_50(oper2[50], oper1[23], g23[50]);
AN2 GA23_51(oper2[51], oper1[23], g23[51]);
AN2 GA23_52(oper2[52], oper1[23], g23[52]);
AN2 GA23_53(oper2[53], oper1[23], g23[53]);
AN2 GA23_54(oper2[54], oper1[23], g23[54]);
AN2 GA23_55(oper2[55], oper1[23], g23[55]);
AN2 GA23_56(oper2[56], oper1[23], g23[56]);
AN2 GA23_57(oper2[57], oper1[23], g23[57]);
AN2 GA23_58(oper2[58], oper1[23], g23[58]);
AN2 GA23_59(oper2[59], oper1[23], g23[59]);
AN2 GA23_60(oper2[60], oper1[23], g23[60]);
AN2 GA23_61(oper2[61], oper1[23], g23[61]);
AN2 GA23_62(oper2[62], oper1[23], g23[62]);
AN2 GA23_63(oper2[63], oper1[23], g23[63]);
AN2 GA22_8(oper2[8], oper1[22], g22[8]);
AN2 GA22_9(oper2[9], oper1[22], g22[9]);
AN2 GA22_10(oper2[10], oper1[22], g22[10]);
AN2 GA22_11(oper2[11], oper1[22], g22[11]);
AN2 GA22_12(oper2[12], oper1[22], g22[12]);
AN2 GA22_13(oper2[13], oper1[22], g22[13]);
AN2 GA22_14(oper2[14], oper1[22], g22[14]);
AN2 GA22_15(oper2[15], oper1[22], g22[15]);
AN2 GA22_16(oper2[16], oper1[22], g22[16]);
AN2 GA22_17(oper2[17], oper1[22], g22[17]);
AN2 GA22_18(oper2[18], oper1[22], g22[18]);
AN2 GA22_19(oper2[19], oper1[22], g22[19]);
AN2 GA22_20(oper2[20], oper1[22], g22[20]);
AN2 GA22_21(oper2[21], oper1[22], g22[21]);
AN2 GA22_22(oper2[22], oper1[22], g22[22]);
AN2 GA22_23(oper2[23], oper1[22], g22[23]);
AN2 GA22_24(oper2[24], oper1[22], g22[24]);
AN2 GA22_25(oper2[25], oper1[22], g22[25]);
AN2 GA22_26(oper2[26], oper1[22], g22[26]);
AN2 GA22_27(oper2[27], oper1[22], g22[27]);
AN2 GA22_28(oper2[28], oper1[22], g22[28]);
AN2 GA22_29(oper2[29], oper1[22], g22[29]);
AN2 GA22_30(oper2[30], oper1[22], g22[30]);
AN2 GA22_31(oper2[31], oper1[22], g22[31]);
AN2 GA22_32(oper2[32], oper1[22], g22[32]);
AN2 GA22_33(oper2[33], oper1[22], g22[33]);
AN2 GA22_34(oper2[34], oper1[22], g22[34]);
AN2 GA22_35(oper2[35], oper1[22], g22[35]);
AN2 GA22_36(oper2[36], oper1[22], g22[36]);
AN2 GA22_37(oper2[37], oper1[22], g22[37]);
AN2 GA22_38(oper2[38], oper1[22], g22[38]);
AN2 GA22_39(oper2[39], oper1[22], g22[39]);
AN2 GA22_40(oper2[40], oper1[22], g22[40]);
AN2 GA22_41(oper2[41], oper1[22], g22[41]);
AN2 GA22_42(oper2[42], oper1[22], g22[42]);
AN2 GA22_43(oper2[43], oper1[22], g22[43]);
AN2 GA22_44(oper2[44], oper1[22], g22[44]);
AN2 GA22_45(oper2[45], oper1[22], g22[45]);
AN2 GA22_46(oper2[46], oper1[22], g22[46]);
AN2 GA22_47(oper2[47], oper1[22], g22[47]);
AN2 GA22_48(oper2[48], oper1[22], g22[48]);
AN2 GA22_49(oper2[49], oper1[22], g22[49]);
AN2 GA22_50(oper2[50], oper1[22], g22[50]);
AN2 GA22_51(oper2[51], oper1[22], g22[51]);
AN2 GA22_52(oper2[52], oper1[22], g22[52]);
AN2 GA22_53(oper2[53], oper1[22], g22[53]);
AN2 GA22_54(oper2[54], oper1[22], g22[54]);
AN2 GA22_55(oper2[55], oper1[22], g22[55]);
AN2 GA22_56(oper2[56], oper1[22], g22[56]);
AN2 GA22_57(oper2[57], oper1[22], g22[57]);
AN2 GA22_58(oper2[58], oper1[22], g22[58]);
AN2 GA22_59(oper2[59], oper1[22], g22[59]);
AN2 GA22_60(oper2[60], oper1[22], g22[60]);
AN2 GA22_61(oper2[61], oper1[22], g22[61]);
AN2 GA22_62(oper2[62], oper1[22], g22[62]);
AN2 GA22_63(oper2[63], oper1[22], g22[63]);
AN2 GA21_8(oper2[8], oper1[21], g21[8]);
AN2 GA21_9(oper2[9], oper1[21], g21[9]);
AN2 GA21_10(oper2[10], oper1[21], g21[10]);
AN2 GA21_11(oper2[11], oper1[21], g21[11]);
AN2 GA21_12(oper2[12], oper1[21], g21[12]);
AN2 GA21_13(oper2[13], oper1[21], g21[13]);
AN2 GA21_14(oper2[14], oper1[21], g21[14]);
AN2 GA21_15(oper2[15], oper1[21], g21[15]);
AN2 GA21_16(oper2[16], oper1[21], g21[16]);
AN2 GA21_17(oper2[17], oper1[21], g21[17]);
AN2 GA21_18(oper2[18], oper1[21], g21[18]);
AN2 GA21_19(oper2[19], oper1[21], g21[19]);
AN2 GA21_20(oper2[20], oper1[21], g21[20]);
AN2 GA21_21(oper2[21], oper1[21], g21[21]);
AN2 GA21_22(oper2[22], oper1[21], g21[22]);
AN2 GA21_23(oper2[23], oper1[21], g21[23]);
AN2 GA21_24(oper2[24], oper1[21], g21[24]);
AN2 GA21_25(oper2[25], oper1[21], g21[25]);
AN2 GA21_26(oper2[26], oper1[21], g21[26]);
AN2 GA21_27(oper2[27], oper1[21], g21[27]);
AN2 GA21_28(oper2[28], oper1[21], g21[28]);
AN2 GA21_29(oper2[29], oper1[21], g21[29]);
AN2 GA21_30(oper2[30], oper1[21], g21[30]);
AN2 GA21_31(oper2[31], oper1[21], g21[31]);
AN2 GA21_32(oper2[32], oper1[21], g21[32]);
AN2 GA21_33(oper2[33], oper1[21], g21[33]);
AN2 GA21_34(oper2[34], oper1[21], g21[34]);
AN2 GA21_35(oper2[35], oper1[21], g21[35]);
AN2 GA21_36(oper2[36], oper1[21], g21[36]);
AN2 GA21_37(oper2[37], oper1[21], g21[37]);
AN2 GA21_38(oper2[38], oper1[21], g21[38]);
AN2 GA21_39(oper2[39], oper1[21], g21[39]);
AN2 GA21_40(oper2[40], oper1[21], g21[40]);
AN2 GA21_41(oper2[41], oper1[21], g21[41]);
AN2 GA21_42(oper2[42], oper1[21], g21[42]);
AN2 GA21_43(oper2[43], oper1[21], g21[43]);
AN2 GA21_44(oper2[44], oper1[21], g21[44]);
AN2 GA21_45(oper2[45], oper1[21], g21[45]);
AN2 GA21_46(oper2[46], oper1[21], g21[46]);
AN2 GA21_47(oper2[47], oper1[21], g21[47]);
AN2 GA21_48(oper2[48], oper1[21], g21[48]);
AN2 GA21_49(oper2[49], oper1[21], g21[49]);
AN2 GA21_50(oper2[50], oper1[21], g21[50]);
AN2 GA21_51(oper2[51], oper1[21], g21[51]);
AN2 GA21_52(oper2[52], oper1[21], g21[52]);
AN2 GA21_53(oper2[53], oper1[21], g21[53]);
AN2 GA21_54(oper2[54], oper1[21], g21[54]);
AN2 GA21_55(oper2[55], oper1[21], g21[55]);
AN2 GA21_56(oper2[56], oper1[21], g21[56]);
AN2 GA21_57(oper2[57], oper1[21], g21[57]);
AN2 GA21_58(oper2[58], oper1[21], g21[58]);
AN2 GA21_59(oper2[59], oper1[21], g21[59]);
AN2 GA21_60(oper2[60], oper1[21], g21[60]);
AN2 GA21_61(oper2[61], oper1[21], g21[61]);
AN2 GA21_62(oper2[62], oper1[21], g21[62]);
AN2 GA21_63(oper2[63], oper1[21], g21[63]);
AN2 GA20_8(oper2[8], oper1[20], g20[8]);
AN2 GA20_9(oper2[9], oper1[20], g20[9]);
AN2 GA20_10(oper2[10], oper1[20], g20[10]);
AN2 GA20_11(oper2[11], oper1[20], g20[11]);
AN2 GA20_12(oper2[12], oper1[20], g20[12]);
AN2 GA20_13(oper2[13], oper1[20], g20[13]);
AN2 GA20_14(oper2[14], oper1[20], g20[14]);
AN2 GA20_15(oper2[15], oper1[20], g20[15]);
AN2 GA20_16(oper2[16], oper1[20], g20[16]);
AN2 GA20_17(oper2[17], oper1[20], g20[17]);
AN2 GA20_18(oper2[18], oper1[20], g20[18]);
AN2 GA20_19(oper2[19], oper1[20], g20[19]);
AN2 GA20_20(oper2[20], oper1[20], g20[20]);
AN2 GA20_21(oper2[21], oper1[20], g20[21]);
AN2 GA20_22(oper2[22], oper1[20], g20[22]);
AN2 GA20_23(oper2[23], oper1[20], g20[23]);
AN2 GA20_24(oper2[24], oper1[20], g20[24]);
AN2 GA20_25(oper2[25], oper1[20], g20[25]);
AN2 GA20_26(oper2[26], oper1[20], g20[26]);
AN2 GA20_27(oper2[27], oper1[20], g20[27]);
AN2 GA20_28(oper2[28], oper1[20], g20[28]);
AN2 GA20_29(oper2[29], oper1[20], g20[29]);
AN2 GA20_30(oper2[30], oper1[20], g20[30]);
AN2 GA20_31(oper2[31], oper1[20], g20[31]);
AN2 GA20_32(oper2[32], oper1[20], g20[32]);
AN2 GA20_33(oper2[33], oper1[20], g20[33]);
AN2 GA20_34(oper2[34], oper1[20], g20[34]);
AN2 GA20_35(oper2[35], oper1[20], g20[35]);
AN2 GA20_36(oper2[36], oper1[20], g20[36]);
AN2 GA20_37(oper2[37], oper1[20], g20[37]);
AN2 GA20_38(oper2[38], oper1[20], g20[38]);
AN2 GA20_39(oper2[39], oper1[20], g20[39]);
AN2 GA20_40(oper2[40], oper1[20], g20[40]);
AN2 GA20_41(oper2[41], oper1[20], g20[41]);
AN2 GA20_42(oper2[42], oper1[20], g20[42]);
AN2 GA20_43(oper2[43], oper1[20], g20[43]);
AN2 GA20_44(oper2[44], oper1[20], g20[44]);
AN2 GA20_45(oper2[45], oper1[20], g20[45]);
AN2 GA20_46(oper2[46], oper1[20], g20[46]);
AN2 GA20_47(oper2[47], oper1[20], g20[47]);
AN2 GA20_48(oper2[48], oper1[20], g20[48]);
AN2 GA20_49(oper2[49], oper1[20], g20[49]);
AN2 GA20_50(oper2[50], oper1[20], g20[50]);
AN2 GA20_51(oper2[51], oper1[20], g20[51]);
AN2 GA20_52(oper2[52], oper1[20], g20[52]);
AN2 GA20_53(oper2[53], oper1[20], g20[53]);
AN2 GA20_54(oper2[54], oper1[20], g20[54]);
AN2 GA20_55(oper2[55], oper1[20], g20[55]);
AN2 GA20_56(oper2[56], oper1[20], g20[56]);
AN2 GA20_57(oper2[57], oper1[20], g20[57]);
AN2 GA20_58(oper2[58], oper1[20], g20[58]);
AN2 GA20_59(oper2[59], oper1[20], g20[59]);
AN2 GA20_60(oper2[60], oper1[20], g20[60]);
AN2 GA20_61(oper2[61], oper1[20], g20[61]);
AN2 GA20_62(oper2[62], oper1[20], g20[62]);
AN2 GA20_63(oper2[63], oper1[20], g20[63]);
AN2 GA19_8(oper2[8], oper1[19], g19[8]);
AN2 GA19_9(oper2[9], oper1[19], g19[9]);
AN2 GA19_10(oper2[10], oper1[19], g19[10]);
AN2 GA19_11(oper2[11], oper1[19], g19[11]);
AN2 GA19_12(oper2[12], oper1[19], g19[12]);
AN2 GA19_13(oper2[13], oper1[19], g19[13]);
AN2 GA19_14(oper2[14], oper1[19], g19[14]);
AN2 GA19_15(oper2[15], oper1[19], g19[15]);
AN2 GA19_16(oper2[16], oper1[19], g19[16]);
AN2 GA19_17(oper2[17], oper1[19], g19[17]);
AN2 GA19_18(oper2[18], oper1[19], g19[18]);
AN2 GA19_19(oper2[19], oper1[19], g19[19]);
AN2 GA19_20(oper2[20], oper1[19], g19[20]);
AN2 GA19_21(oper2[21], oper1[19], g19[21]);
AN2 GA19_22(oper2[22], oper1[19], g19[22]);
AN2 GA19_23(oper2[23], oper1[19], g19[23]);
AN2 GA19_24(oper2[24], oper1[19], g19[24]);
AN2 GA19_25(oper2[25], oper1[19], g19[25]);
AN2 GA19_26(oper2[26], oper1[19], g19[26]);
AN2 GA19_27(oper2[27], oper1[19], g19[27]);
AN2 GA19_28(oper2[28], oper1[19], g19[28]);
AN2 GA19_29(oper2[29], oper1[19], g19[29]);
AN2 GA19_30(oper2[30], oper1[19], g19[30]);
AN2 GA19_31(oper2[31], oper1[19], g19[31]);
AN2 GA19_32(oper2[32], oper1[19], g19[32]);
AN2 GA19_33(oper2[33], oper1[19], g19[33]);
AN2 GA19_34(oper2[34], oper1[19], g19[34]);
AN2 GA19_35(oper2[35], oper1[19], g19[35]);
AN2 GA19_36(oper2[36], oper1[19], g19[36]);
AN2 GA19_37(oper2[37], oper1[19], g19[37]);
AN2 GA19_38(oper2[38], oper1[19], g19[38]);
AN2 GA19_39(oper2[39], oper1[19], g19[39]);
AN2 GA19_40(oper2[40], oper1[19], g19[40]);
AN2 GA19_41(oper2[41], oper1[19], g19[41]);
AN2 GA19_42(oper2[42], oper1[19], g19[42]);
AN2 GA19_43(oper2[43], oper1[19], g19[43]);
AN2 GA19_44(oper2[44], oper1[19], g19[44]);
AN2 GA19_45(oper2[45], oper1[19], g19[45]);
AN2 GA19_46(oper2[46], oper1[19], g19[46]);
AN2 GA19_47(oper2[47], oper1[19], g19[47]);
AN2 GA19_48(oper2[48], oper1[19], g19[48]);
AN2 GA19_49(oper2[49], oper1[19], g19[49]);
AN2 GA19_50(oper2[50], oper1[19], g19[50]);
AN2 GA19_51(oper2[51], oper1[19], g19[51]);
AN2 GA19_52(oper2[52], oper1[19], g19[52]);
AN2 GA19_53(oper2[53], oper1[19], g19[53]);
AN2 GA19_54(oper2[54], oper1[19], g19[54]);
AN2 GA19_55(oper2[55], oper1[19], g19[55]);
AN2 GA19_56(oper2[56], oper1[19], g19[56]);
AN2 GA19_57(oper2[57], oper1[19], g19[57]);
AN2 GA19_58(oper2[58], oper1[19], g19[58]);
AN2 GA19_59(oper2[59], oper1[19], g19[59]);
AN2 GA19_60(oper2[60], oper1[19], g19[60]);
AN2 GA19_61(oper2[61], oper1[19], g19[61]);
AN2 GA19_62(oper2[62], oper1[19], g19[62]);
AN2 GA19_63(oper2[63], oper1[19], g19[63]);
AN2 GA18_8(oper2[8], oper1[18], g18[8]);
AN2 GA18_9(oper2[9], oper1[18], g18[9]);
AN2 GA18_10(oper2[10], oper1[18], g18[10]);
AN2 GA18_11(oper2[11], oper1[18], g18[11]);
AN2 GA18_12(oper2[12], oper1[18], g18[12]);
AN2 GA18_13(oper2[13], oper1[18], g18[13]);
AN2 GA18_14(oper2[14], oper1[18], g18[14]);
AN2 GA18_15(oper2[15], oper1[18], g18[15]);
AN2 GA18_16(oper2[16], oper1[18], g18[16]);
AN2 GA18_17(oper2[17], oper1[18], g18[17]);
AN2 GA18_18(oper2[18], oper1[18], g18[18]);
AN2 GA18_19(oper2[19], oper1[18], g18[19]);
AN2 GA18_20(oper2[20], oper1[18], g18[20]);
AN2 GA18_21(oper2[21], oper1[18], g18[21]);
AN2 GA18_22(oper2[22], oper1[18], g18[22]);
AN2 GA18_23(oper2[23], oper1[18], g18[23]);
AN2 GA18_24(oper2[24], oper1[18], g18[24]);
AN2 GA18_25(oper2[25], oper1[18], g18[25]);
AN2 GA18_26(oper2[26], oper1[18], g18[26]);
AN2 GA18_27(oper2[27], oper1[18], g18[27]);
AN2 GA18_28(oper2[28], oper1[18], g18[28]);
AN2 GA18_29(oper2[29], oper1[18], g18[29]);
AN2 GA18_30(oper2[30], oper1[18], g18[30]);
AN2 GA18_31(oper2[31], oper1[18], g18[31]);
AN2 GA18_32(oper2[32], oper1[18], g18[32]);
AN2 GA18_33(oper2[33], oper1[18], g18[33]);
AN2 GA18_34(oper2[34], oper1[18], g18[34]);
AN2 GA18_35(oper2[35], oper1[18], g18[35]);
AN2 GA18_36(oper2[36], oper1[18], g18[36]);
AN2 GA18_37(oper2[37], oper1[18], g18[37]);
AN2 GA18_38(oper2[38], oper1[18], g18[38]);
AN2 GA18_39(oper2[39], oper1[18], g18[39]);
AN2 GA18_40(oper2[40], oper1[18], g18[40]);
AN2 GA18_41(oper2[41], oper1[18], g18[41]);
AN2 GA18_42(oper2[42], oper1[18], g18[42]);
AN2 GA18_43(oper2[43], oper1[18], g18[43]);
AN2 GA18_44(oper2[44], oper1[18], g18[44]);
AN2 GA18_45(oper2[45], oper1[18], g18[45]);
AN2 GA18_46(oper2[46], oper1[18], g18[46]);
AN2 GA18_47(oper2[47], oper1[18], g18[47]);
AN2 GA18_48(oper2[48], oper1[18], g18[48]);
AN2 GA18_49(oper2[49], oper1[18], g18[49]);
AN2 GA18_50(oper2[50], oper1[18], g18[50]);
AN2 GA18_51(oper2[51], oper1[18], g18[51]);
AN2 GA18_52(oper2[52], oper1[18], g18[52]);
AN2 GA18_53(oper2[53], oper1[18], g18[53]);
AN2 GA18_54(oper2[54], oper1[18], g18[54]);
AN2 GA18_55(oper2[55], oper1[18], g18[55]);
AN2 GA18_56(oper2[56], oper1[18], g18[56]);
AN2 GA18_57(oper2[57], oper1[18], g18[57]);
AN2 GA18_58(oper2[58], oper1[18], g18[58]);
AN2 GA18_59(oper2[59], oper1[18], g18[59]);
AN2 GA18_60(oper2[60], oper1[18], g18[60]);
AN2 GA18_61(oper2[61], oper1[18], g18[61]);
AN2 GA18_62(oper2[62], oper1[18], g18[62]);
AN2 GA18_63(oper2[63], oper1[18], g18[63]);
AN2 GA17_8(oper2[8], oper1[17], g17[8]);
AN2 GA17_9(oper2[9], oper1[17], g17[9]);
AN2 GA17_10(oper2[10], oper1[17], g17[10]);
AN2 GA17_11(oper2[11], oper1[17], g17[11]);
AN2 GA17_12(oper2[12], oper1[17], g17[12]);
AN2 GA17_13(oper2[13], oper1[17], g17[13]);
AN2 GA17_14(oper2[14], oper1[17], g17[14]);
AN2 GA17_15(oper2[15], oper1[17], g17[15]);
AN2 GA17_16(oper2[16], oper1[17], g17[16]);
AN2 GA17_17(oper2[17], oper1[17], g17[17]);
AN2 GA17_18(oper2[18], oper1[17], g17[18]);
AN2 GA17_19(oper2[19], oper1[17], g17[19]);
AN2 GA17_20(oper2[20], oper1[17], g17[20]);
AN2 GA17_21(oper2[21], oper1[17], g17[21]);
AN2 GA17_22(oper2[22], oper1[17], g17[22]);
AN2 GA17_23(oper2[23], oper1[17], g17[23]);
AN2 GA17_24(oper2[24], oper1[17], g17[24]);
AN2 GA17_25(oper2[25], oper1[17], g17[25]);
AN2 GA17_26(oper2[26], oper1[17], g17[26]);
AN2 GA17_27(oper2[27], oper1[17], g17[27]);
AN2 GA17_28(oper2[28], oper1[17], g17[28]);
AN2 GA17_29(oper2[29], oper1[17], g17[29]);
AN2 GA17_30(oper2[30], oper1[17], g17[30]);
AN2 GA17_31(oper2[31], oper1[17], g17[31]);
AN2 GA17_32(oper2[32], oper1[17], g17[32]);
AN2 GA17_33(oper2[33], oper1[17], g17[33]);
AN2 GA17_34(oper2[34], oper1[17], g17[34]);
AN2 GA17_35(oper2[35], oper1[17], g17[35]);
AN2 GA17_36(oper2[36], oper1[17], g17[36]);
AN2 GA17_37(oper2[37], oper1[17], g17[37]);
AN2 GA17_38(oper2[38], oper1[17], g17[38]);
AN2 GA17_39(oper2[39], oper1[17], g17[39]);
AN2 GA17_40(oper2[40], oper1[17], g17[40]);
AN2 GA17_41(oper2[41], oper1[17], g17[41]);
AN2 GA17_42(oper2[42], oper1[17], g17[42]);
AN2 GA17_43(oper2[43], oper1[17], g17[43]);
AN2 GA17_44(oper2[44], oper1[17], g17[44]);
AN2 GA17_45(oper2[45], oper1[17], g17[45]);
AN2 GA17_46(oper2[46], oper1[17], g17[46]);
AN2 GA17_47(oper2[47], oper1[17], g17[47]);
AN2 GA17_48(oper2[48], oper1[17], g17[48]);
AN2 GA17_49(oper2[49], oper1[17], g17[49]);
AN2 GA17_50(oper2[50], oper1[17], g17[50]);
AN2 GA17_51(oper2[51], oper1[17], g17[51]);
AN2 GA17_52(oper2[52], oper1[17], g17[52]);
AN2 GA17_53(oper2[53], oper1[17], g17[53]);
AN2 GA17_54(oper2[54], oper1[17], g17[54]);
AN2 GA17_55(oper2[55], oper1[17], g17[55]);
AN2 GA17_56(oper2[56], oper1[17], g17[56]);
AN2 GA17_57(oper2[57], oper1[17], g17[57]);
AN2 GA17_58(oper2[58], oper1[17], g17[58]);
AN2 GA17_59(oper2[59], oper1[17], g17[59]);
AN2 GA17_60(oper2[60], oper1[17], g17[60]);
AN2 GA17_61(oper2[61], oper1[17], g17[61]);
AN2 GA17_62(oper2[62], oper1[17], g17[62]);
AN2 GA17_63(oper2[63], oper1[17], g17[63]);
AN2 GA16_8(oper2[8], oper1[16], g16[8]);
AN2 GA16_9(oper2[9], oper1[16], g16[9]);
AN2 GA16_10(oper2[10], oper1[16], g16[10]);
AN2 GA16_11(oper2[11], oper1[16], g16[11]);
AN2 GA16_12(oper2[12], oper1[16], g16[12]);
AN2 GA16_13(oper2[13], oper1[16], g16[13]);
AN2 GA16_14(oper2[14], oper1[16], g16[14]);
AN2 GA16_15(oper2[15], oper1[16], g16[15]);
AN2 GA16_16(oper2[16], oper1[16], g16[16]);
AN2 GA16_17(oper2[17], oper1[16], g16[17]);
AN2 GA16_18(oper2[18], oper1[16], g16[18]);
AN2 GA16_19(oper2[19], oper1[16], g16[19]);
AN2 GA16_20(oper2[20], oper1[16], g16[20]);
AN2 GA16_21(oper2[21], oper1[16], g16[21]);
AN2 GA16_22(oper2[22], oper1[16], g16[22]);
AN2 GA16_23(oper2[23], oper1[16], g16[23]);
AN2 GA16_24(oper2[24], oper1[16], g16[24]);
AN2 GA16_25(oper2[25], oper1[16], g16[25]);
AN2 GA16_26(oper2[26], oper1[16], g16[26]);
AN2 GA16_27(oper2[27], oper1[16], g16[27]);
AN2 GA16_28(oper2[28], oper1[16], g16[28]);
AN2 GA16_29(oper2[29], oper1[16], g16[29]);
AN2 GA16_30(oper2[30], oper1[16], g16[30]);
AN2 GA16_31(oper2[31], oper1[16], g16[31]);
AN2 GA16_32(oper2[32], oper1[16], g16[32]);
AN2 GA16_33(oper2[33], oper1[16], g16[33]);
AN2 GA16_34(oper2[34], oper1[16], g16[34]);
AN2 GA16_35(oper2[35], oper1[16], g16[35]);
AN2 GA16_36(oper2[36], oper1[16], g16[36]);
AN2 GA16_37(oper2[37], oper1[16], g16[37]);
AN2 GA16_38(oper2[38], oper1[16], g16[38]);
AN2 GA16_39(oper2[39], oper1[16], g16[39]);
AN2 GA16_40(oper2[40], oper1[16], g16[40]);
AN2 GA16_41(oper2[41], oper1[16], g16[41]);
AN2 GA16_42(oper2[42], oper1[16], g16[42]);
AN2 GA16_43(oper2[43], oper1[16], g16[43]);
AN2 GA16_44(oper2[44], oper1[16], g16[44]);
AN2 GA16_45(oper2[45], oper1[16], g16[45]);
AN2 GA16_46(oper2[46], oper1[16], g16[46]);
AN2 GA16_47(oper2[47], oper1[16], g16[47]);
AN2 GA16_48(oper2[48], oper1[16], g16[48]);
AN2 GA16_49(oper2[49], oper1[16], g16[49]);
AN2 GA16_50(oper2[50], oper1[16], g16[50]);
AN2 GA16_51(oper2[51], oper1[16], g16[51]);
AN2 GA16_52(oper2[52], oper1[16], g16[52]);
AN2 GA16_53(oper2[53], oper1[16], g16[53]);
AN2 GA16_54(oper2[54], oper1[16], g16[54]);
AN2 GA16_55(oper2[55], oper1[16], g16[55]);
AN2 GA16_56(oper2[56], oper1[16], g16[56]);
AN2 GA16_57(oper2[57], oper1[16], g16[57]);
AN2 GA16_58(oper2[58], oper1[16], g16[58]);
AN2 GA16_59(oper2[59], oper1[16], g16[59]);
AN2 GA16_60(oper2[60], oper1[16], g16[60]);
AN2 GA16_61(oper2[61], oper1[16], g16[61]);
AN2 GA16_62(oper2[62], oper1[16], g16[62]);
AN2 GA16_63(oper2[63], oper1[16], g16[63]);
AN2 GA15_8(oper2[8], oper1[15], g15[8]);
AN2 GA15_9(oper2[9], oper1[15], g15[9]);
AN2 GA15_10(oper2[10], oper1[15], g15[10]);
AN2 GA15_11(oper2[11], oper1[15], g15[11]);
AN2 GA15_12(oper2[12], oper1[15], g15[12]);
AN2 GA15_13(oper2[13], oper1[15], g15[13]);
AN2 GA15_14(oper2[14], oper1[15], g15[14]);
AN2 GA15_15(oper2[15], oper1[15], g15[15]);
AN2 GA15_16(oper2[16], oper1[15], g15[16]);
AN2 GA15_17(oper2[17], oper1[15], g15[17]);
AN2 GA15_18(oper2[18], oper1[15], g15[18]);
AN2 GA15_19(oper2[19], oper1[15], g15[19]);
AN2 GA15_20(oper2[20], oper1[15], g15[20]);
AN2 GA15_21(oper2[21], oper1[15], g15[21]);
AN2 GA15_22(oper2[22], oper1[15], g15[22]);
AN2 GA15_23(oper2[23], oper1[15], g15[23]);
AN2 GA15_24(oper2[24], oper1[15], g15[24]);
AN2 GA15_25(oper2[25], oper1[15], g15[25]);
AN2 GA15_26(oper2[26], oper1[15], g15[26]);
AN2 GA15_27(oper2[27], oper1[15], g15[27]);
AN2 GA15_28(oper2[28], oper1[15], g15[28]);
AN2 GA15_29(oper2[29], oper1[15], g15[29]);
AN2 GA15_30(oper2[30], oper1[15], g15[30]);
AN2 GA15_31(oper2[31], oper1[15], g15[31]);
AN2 GA15_32(oper2[32], oper1[15], g15[32]);
AN2 GA15_33(oper2[33], oper1[15], g15[33]);
AN2 GA15_34(oper2[34], oper1[15], g15[34]);
AN2 GA15_35(oper2[35], oper1[15], g15[35]);
AN2 GA15_36(oper2[36], oper1[15], g15[36]);
AN2 GA15_37(oper2[37], oper1[15], g15[37]);
AN2 GA15_38(oper2[38], oper1[15], g15[38]);
AN2 GA15_39(oper2[39], oper1[15], g15[39]);
AN2 GA15_40(oper2[40], oper1[15], g15[40]);
AN2 GA15_41(oper2[41], oper1[15], g15[41]);
AN2 GA15_42(oper2[42], oper1[15], g15[42]);
AN2 GA15_43(oper2[43], oper1[15], g15[43]);
AN2 GA15_44(oper2[44], oper1[15], g15[44]);
AN2 GA15_45(oper2[45], oper1[15], g15[45]);
AN2 GA15_46(oper2[46], oper1[15], g15[46]);
AN2 GA15_47(oper2[47], oper1[15], g15[47]);
AN2 GA15_48(oper2[48], oper1[15], g15[48]);
AN2 GA15_49(oper2[49], oper1[15], g15[49]);
AN2 GA15_50(oper2[50], oper1[15], g15[50]);
AN2 GA15_51(oper2[51], oper1[15], g15[51]);
AN2 GA15_52(oper2[52], oper1[15], g15[52]);
AN2 GA15_53(oper2[53], oper1[15], g15[53]);
AN2 GA15_54(oper2[54], oper1[15], g15[54]);
AN2 GA15_55(oper2[55], oper1[15], g15[55]);
AN2 GA15_56(oper2[56], oper1[15], g15[56]);
AN2 GA15_57(oper2[57], oper1[15], g15[57]);
AN2 GA15_58(oper2[58], oper1[15], g15[58]);
AN2 GA15_59(oper2[59], oper1[15], g15[59]);
AN2 GA15_60(oper2[60], oper1[15], g15[60]);
AN2 GA15_61(oper2[61], oper1[15], g15[61]);
AN2 GA15_62(oper2[62], oper1[15], g15[62]);
AN2 GA15_63(oper2[63], oper1[15], g15[63]);
AN2 GA14_8(oper2[8], oper1[14], g14[8]);
AN2 GA14_9(oper2[9], oper1[14], g14[9]);
AN2 GA14_10(oper2[10], oper1[14], g14[10]);
AN2 GA14_11(oper2[11], oper1[14], g14[11]);
AN2 GA14_12(oper2[12], oper1[14], g14[12]);
AN2 GA14_13(oper2[13], oper1[14], g14[13]);
AN2 GA14_14(oper2[14], oper1[14], g14[14]);
AN2 GA14_15(oper2[15], oper1[14], g14[15]);
AN2 GA14_16(oper2[16], oper1[14], g14[16]);
AN2 GA14_17(oper2[17], oper1[14], g14[17]);
AN2 GA14_18(oper2[18], oper1[14], g14[18]);
AN2 GA14_19(oper2[19], oper1[14], g14[19]);
AN2 GA14_20(oper2[20], oper1[14], g14[20]);
AN2 GA14_21(oper2[21], oper1[14], g14[21]);
AN2 GA14_22(oper2[22], oper1[14], g14[22]);
AN2 GA14_23(oper2[23], oper1[14], g14[23]);
AN2 GA14_24(oper2[24], oper1[14], g14[24]);
AN2 GA14_25(oper2[25], oper1[14], g14[25]);
AN2 GA14_26(oper2[26], oper1[14], g14[26]);
AN2 GA14_27(oper2[27], oper1[14], g14[27]);
AN2 GA14_28(oper2[28], oper1[14], g14[28]);
AN2 GA14_29(oper2[29], oper1[14], g14[29]);
AN2 GA14_30(oper2[30], oper1[14], g14[30]);
AN2 GA14_31(oper2[31], oper1[14], g14[31]);
AN2 GA14_32(oper2[32], oper1[14], g14[32]);
AN2 GA14_33(oper2[33], oper1[14], g14[33]);
AN2 GA14_34(oper2[34], oper1[14], g14[34]);
AN2 GA14_35(oper2[35], oper1[14], g14[35]);
AN2 GA14_36(oper2[36], oper1[14], g14[36]);
AN2 GA14_37(oper2[37], oper1[14], g14[37]);
AN2 GA14_38(oper2[38], oper1[14], g14[38]);
AN2 GA14_39(oper2[39], oper1[14], g14[39]);
AN2 GA14_40(oper2[40], oper1[14], g14[40]);
AN2 GA14_41(oper2[41], oper1[14], g14[41]);
AN2 GA14_42(oper2[42], oper1[14], g14[42]);
AN2 GA14_43(oper2[43], oper1[14], g14[43]);
AN2 GA14_44(oper2[44], oper1[14], g14[44]);
AN2 GA14_45(oper2[45], oper1[14], g14[45]);
AN2 GA14_46(oper2[46], oper1[14], g14[46]);
AN2 GA14_47(oper2[47], oper1[14], g14[47]);
AN2 GA14_48(oper2[48], oper1[14], g14[48]);
AN2 GA14_49(oper2[49], oper1[14], g14[49]);
AN2 GA14_50(oper2[50], oper1[14], g14[50]);
AN2 GA14_51(oper2[51], oper1[14], g14[51]);
AN2 GA14_52(oper2[52], oper1[14], g14[52]);
AN2 GA14_53(oper2[53], oper1[14], g14[53]);
AN2 GA14_54(oper2[54], oper1[14], g14[54]);
AN2 GA14_55(oper2[55], oper1[14], g14[55]);
AN2 GA14_56(oper2[56], oper1[14], g14[56]);
AN2 GA14_57(oper2[57], oper1[14], g14[57]);
AN2 GA14_58(oper2[58], oper1[14], g14[58]);
AN2 GA14_59(oper2[59], oper1[14], g14[59]);
AN2 GA14_60(oper2[60], oper1[14], g14[60]);
AN2 GA14_61(oper2[61], oper1[14], g14[61]);
AN2 GA14_62(oper2[62], oper1[14], g14[62]);
AN2 GA14_63(oper2[63], oper1[14], g14[63]);
AN2 GA13_8(oper2[8], oper1[13], g13[8]);
AN2 GA13_9(oper2[9], oper1[13], g13[9]);
AN2 GA13_10(oper2[10], oper1[13], g13[10]);
AN2 GA13_11(oper2[11], oper1[13], g13[11]);
AN2 GA13_12(oper2[12], oper1[13], g13[12]);
AN2 GA13_13(oper2[13], oper1[13], g13[13]);
AN2 GA13_14(oper2[14], oper1[13], g13[14]);
AN2 GA13_15(oper2[15], oper1[13], g13[15]);
AN2 GA13_16(oper2[16], oper1[13], g13[16]);
AN2 GA13_17(oper2[17], oper1[13], g13[17]);
AN2 GA13_18(oper2[18], oper1[13], g13[18]);
AN2 GA13_19(oper2[19], oper1[13], g13[19]);
AN2 GA13_20(oper2[20], oper1[13], g13[20]);
AN2 GA13_21(oper2[21], oper1[13], g13[21]);
AN2 GA13_22(oper2[22], oper1[13], g13[22]);
AN2 GA13_23(oper2[23], oper1[13], g13[23]);
AN2 GA13_24(oper2[24], oper1[13], g13[24]);
AN2 GA13_25(oper2[25], oper1[13], g13[25]);
AN2 GA13_26(oper2[26], oper1[13], g13[26]);
AN2 GA13_27(oper2[27], oper1[13], g13[27]);
AN2 GA13_28(oper2[28], oper1[13], g13[28]);
AN2 GA13_29(oper2[29], oper1[13], g13[29]);
AN2 GA13_30(oper2[30], oper1[13], g13[30]);
AN2 GA13_31(oper2[31], oper1[13], g13[31]);
AN2 GA13_32(oper2[32], oper1[13], g13[32]);
AN2 GA13_33(oper2[33], oper1[13], g13[33]);
AN2 GA13_34(oper2[34], oper1[13], g13[34]);
AN2 GA13_35(oper2[35], oper1[13], g13[35]);
AN2 GA13_36(oper2[36], oper1[13], g13[36]);
AN2 GA13_37(oper2[37], oper1[13], g13[37]);
AN2 GA13_38(oper2[38], oper1[13], g13[38]);
AN2 GA13_39(oper2[39], oper1[13], g13[39]);
AN2 GA13_40(oper2[40], oper1[13], g13[40]);
AN2 GA13_41(oper2[41], oper1[13], g13[41]);
AN2 GA13_42(oper2[42], oper1[13], g13[42]);
AN2 GA13_43(oper2[43], oper1[13], g13[43]);
AN2 GA13_44(oper2[44], oper1[13], g13[44]);
AN2 GA13_45(oper2[45], oper1[13], g13[45]);
AN2 GA13_46(oper2[46], oper1[13], g13[46]);
AN2 GA13_47(oper2[47], oper1[13], g13[47]);
AN2 GA13_48(oper2[48], oper1[13], g13[48]);
AN2 GA13_49(oper2[49], oper1[13], g13[49]);
AN2 GA13_50(oper2[50], oper1[13], g13[50]);
AN2 GA13_51(oper2[51], oper1[13], g13[51]);
AN2 GA13_52(oper2[52], oper1[13], g13[52]);
AN2 GA13_53(oper2[53], oper1[13], g13[53]);
AN2 GA13_54(oper2[54], oper1[13], g13[54]);
AN2 GA13_55(oper2[55], oper1[13], g13[55]);
AN2 GA13_56(oper2[56], oper1[13], g13[56]);
AN2 GA13_57(oper2[57], oper1[13], g13[57]);
AN2 GA13_58(oper2[58], oper1[13], g13[58]);
AN2 GA13_59(oper2[59], oper1[13], g13[59]);
AN2 GA13_60(oper2[60], oper1[13], g13[60]);
AN2 GA13_61(oper2[61], oper1[13], g13[61]);
AN2 GA13_62(oper2[62], oper1[13], g13[62]);
AN2 GA13_63(oper2[63], oper1[13], g13[63]);
AN2 GA12_8(oper2[8], oper1[12], g12[8]);
AN2 GA12_9(oper2[9], oper1[12], g12[9]);
AN2 GA12_10(oper2[10], oper1[12], g12[10]);
AN2 GA12_11(oper2[11], oper1[12], g12[11]);
AN2 GA12_12(oper2[12], oper1[12], g12[12]);
AN2 GA12_13(oper2[13], oper1[12], g12[13]);
AN2 GA12_14(oper2[14], oper1[12], g12[14]);
AN2 GA12_15(oper2[15], oper1[12], g12[15]);
AN2 GA12_16(oper2[16], oper1[12], g12[16]);
AN2 GA12_17(oper2[17], oper1[12], g12[17]);
AN2 GA12_18(oper2[18], oper1[12], g12[18]);
AN2 GA12_19(oper2[19], oper1[12], g12[19]);
AN2 GA12_20(oper2[20], oper1[12], g12[20]);
AN2 GA12_21(oper2[21], oper1[12], g12[21]);
AN2 GA12_22(oper2[22], oper1[12], g12[22]);
AN2 GA12_23(oper2[23], oper1[12], g12[23]);
AN2 GA12_24(oper2[24], oper1[12], g12[24]);
AN2 GA12_25(oper2[25], oper1[12], g12[25]);
AN2 GA12_26(oper2[26], oper1[12], g12[26]);
AN2 GA12_27(oper2[27], oper1[12], g12[27]);
AN2 GA12_28(oper2[28], oper1[12], g12[28]);
AN2 GA12_29(oper2[29], oper1[12], g12[29]);
AN2 GA12_30(oper2[30], oper1[12], g12[30]);
AN2 GA12_31(oper2[31], oper1[12], g12[31]);
AN2 GA12_32(oper2[32], oper1[12], g12[32]);
AN2 GA12_33(oper2[33], oper1[12], g12[33]);
AN2 GA12_34(oper2[34], oper1[12], g12[34]);
AN2 GA12_35(oper2[35], oper1[12], g12[35]);
AN2 GA12_36(oper2[36], oper1[12], g12[36]);
AN2 GA12_37(oper2[37], oper1[12], g12[37]);
AN2 GA12_38(oper2[38], oper1[12], g12[38]);
AN2 GA12_39(oper2[39], oper1[12], g12[39]);
AN2 GA12_40(oper2[40], oper1[12], g12[40]);
AN2 GA12_41(oper2[41], oper1[12], g12[41]);
AN2 GA12_42(oper2[42], oper1[12], g12[42]);
AN2 GA12_43(oper2[43], oper1[12], g12[43]);
AN2 GA12_44(oper2[44], oper1[12], g12[44]);
AN2 GA12_45(oper2[45], oper1[12], g12[45]);
AN2 GA12_46(oper2[46], oper1[12], g12[46]);
AN2 GA12_47(oper2[47], oper1[12], g12[47]);
AN2 GA12_48(oper2[48], oper1[12], g12[48]);
AN2 GA12_49(oper2[49], oper1[12], g12[49]);
AN2 GA12_50(oper2[50], oper1[12], g12[50]);
AN2 GA12_51(oper2[51], oper1[12], g12[51]);
AN2 GA12_52(oper2[52], oper1[12], g12[52]);
AN2 GA12_53(oper2[53], oper1[12], g12[53]);
AN2 GA12_54(oper2[54], oper1[12], g12[54]);
AN2 GA12_55(oper2[55], oper1[12], g12[55]);
AN2 GA12_56(oper2[56], oper1[12], g12[56]);
AN2 GA12_57(oper2[57], oper1[12], g12[57]);
AN2 GA12_58(oper2[58], oper1[12], g12[58]);
AN2 GA12_59(oper2[59], oper1[12], g12[59]);
AN2 GA12_60(oper2[60], oper1[12], g12[60]);
AN2 GA12_61(oper2[61], oper1[12], g12[61]);
AN2 GA12_62(oper2[62], oper1[12], g12[62]);
AN2 GA12_63(oper2[63], oper1[12], g12[63]);
AN2 GA11_8(oper2[8], oper1[11], g11[8]);
AN2 GA11_9(oper2[9], oper1[11], g11[9]);
AN2 GA11_10(oper2[10], oper1[11], g11[10]);
AN2 GA11_11(oper2[11], oper1[11], g11[11]);
AN2 GA11_12(oper2[12], oper1[11], g11[12]);
AN2 GA11_13(oper2[13], oper1[11], g11[13]);
AN2 GA11_14(oper2[14], oper1[11], g11[14]);
AN2 GA11_15(oper2[15], oper1[11], g11[15]);
AN2 GA11_16(oper2[16], oper1[11], g11[16]);
AN2 GA11_17(oper2[17], oper1[11], g11[17]);
AN2 GA11_18(oper2[18], oper1[11], g11[18]);
AN2 GA11_19(oper2[19], oper1[11], g11[19]);
AN2 GA11_20(oper2[20], oper1[11], g11[20]);
AN2 GA11_21(oper2[21], oper1[11], g11[21]);
AN2 GA11_22(oper2[22], oper1[11], g11[22]);
AN2 GA11_23(oper2[23], oper1[11], g11[23]);
AN2 GA11_24(oper2[24], oper1[11], g11[24]);
AN2 GA11_25(oper2[25], oper1[11], g11[25]);
AN2 GA11_26(oper2[26], oper1[11], g11[26]);
AN2 GA11_27(oper2[27], oper1[11], g11[27]);
AN2 GA11_28(oper2[28], oper1[11], g11[28]);
AN2 GA11_29(oper2[29], oper1[11], g11[29]);
AN2 GA11_30(oper2[30], oper1[11], g11[30]);
AN2 GA11_31(oper2[31], oper1[11], g11[31]);
AN2 GA11_32(oper2[32], oper1[11], g11[32]);
AN2 GA11_33(oper2[33], oper1[11], g11[33]);
AN2 GA11_34(oper2[34], oper1[11], g11[34]);
AN2 GA11_35(oper2[35], oper1[11], g11[35]);
AN2 GA11_36(oper2[36], oper1[11], g11[36]);
AN2 GA11_37(oper2[37], oper1[11], g11[37]);
AN2 GA11_38(oper2[38], oper1[11], g11[38]);
AN2 GA11_39(oper2[39], oper1[11], g11[39]);
AN2 GA11_40(oper2[40], oper1[11], g11[40]);
AN2 GA11_41(oper2[41], oper1[11], g11[41]);
AN2 GA11_42(oper2[42], oper1[11], g11[42]);
AN2 GA11_43(oper2[43], oper1[11], g11[43]);
AN2 GA11_44(oper2[44], oper1[11], g11[44]);
AN2 GA11_45(oper2[45], oper1[11], g11[45]);
AN2 GA11_46(oper2[46], oper1[11], g11[46]);
AN2 GA11_47(oper2[47], oper1[11], g11[47]);
AN2 GA11_48(oper2[48], oper1[11], g11[48]);
AN2 GA11_49(oper2[49], oper1[11], g11[49]);
AN2 GA11_50(oper2[50], oper1[11], g11[50]);
AN2 GA11_51(oper2[51], oper1[11], g11[51]);
AN2 GA11_52(oper2[52], oper1[11], g11[52]);
AN2 GA11_53(oper2[53], oper1[11], g11[53]);
AN2 GA11_54(oper2[54], oper1[11], g11[54]);
AN2 GA11_55(oper2[55], oper1[11], g11[55]);
AN2 GA11_56(oper2[56], oper1[11], g11[56]);
AN2 GA11_57(oper2[57], oper1[11], g11[57]);
AN2 GA11_58(oper2[58], oper1[11], g11[58]);
AN2 GA11_59(oper2[59], oper1[11], g11[59]);
AN2 GA11_60(oper2[60], oper1[11], g11[60]);
AN2 GA11_61(oper2[61], oper1[11], g11[61]);
AN2 GA11_62(oper2[62], oper1[11], g11[62]);
AN2 GA11_63(oper2[63], oper1[11], g11[63]);
AN2 GA10_8(oper2[8], oper1[10], g10[8]);
AN2 GA10_9(oper2[9], oper1[10], g10[9]);
AN2 GA10_10(oper2[10], oper1[10], g10[10]);
AN2 GA10_11(oper2[11], oper1[10], g10[11]);
AN2 GA10_12(oper2[12], oper1[10], g10[12]);
AN2 GA10_13(oper2[13], oper1[10], g10[13]);
AN2 GA10_14(oper2[14], oper1[10], g10[14]);
AN2 GA10_15(oper2[15], oper1[10], g10[15]);
AN2 GA10_16(oper2[16], oper1[10], g10[16]);
AN2 GA10_17(oper2[17], oper1[10], g10[17]);
AN2 GA10_18(oper2[18], oper1[10], g10[18]);
AN2 GA10_19(oper2[19], oper1[10], g10[19]);
AN2 GA10_20(oper2[20], oper1[10], g10[20]);
AN2 GA10_21(oper2[21], oper1[10], g10[21]);
AN2 GA10_22(oper2[22], oper1[10], g10[22]);
AN2 GA10_23(oper2[23], oper1[10], g10[23]);
AN2 GA10_24(oper2[24], oper1[10], g10[24]);
AN2 GA10_25(oper2[25], oper1[10], g10[25]);
AN2 GA10_26(oper2[26], oper1[10], g10[26]);
AN2 GA10_27(oper2[27], oper1[10], g10[27]);
AN2 GA10_28(oper2[28], oper1[10], g10[28]);
AN2 GA10_29(oper2[29], oper1[10], g10[29]);
AN2 GA10_30(oper2[30], oper1[10], g10[30]);
AN2 GA10_31(oper2[31], oper1[10], g10[31]);
AN2 GA10_32(oper2[32], oper1[10], g10[32]);
AN2 GA10_33(oper2[33], oper1[10], g10[33]);
AN2 GA10_34(oper2[34], oper1[10], g10[34]);
AN2 GA10_35(oper2[35], oper1[10], g10[35]);
AN2 GA10_36(oper2[36], oper1[10], g10[36]);
AN2 GA10_37(oper2[37], oper1[10], g10[37]);
AN2 GA10_38(oper2[38], oper1[10], g10[38]);
AN2 GA10_39(oper2[39], oper1[10], g10[39]);
AN2 GA10_40(oper2[40], oper1[10], g10[40]);
AN2 GA10_41(oper2[41], oper1[10], g10[41]);
AN2 GA10_42(oper2[42], oper1[10], g10[42]);
AN2 GA10_43(oper2[43], oper1[10], g10[43]);
AN2 GA10_44(oper2[44], oper1[10], g10[44]);
AN2 GA10_45(oper2[45], oper1[10], g10[45]);
AN2 GA10_46(oper2[46], oper1[10], g10[46]);
AN2 GA10_47(oper2[47], oper1[10], g10[47]);
AN2 GA10_48(oper2[48], oper1[10], g10[48]);
AN2 GA10_49(oper2[49], oper1[10], g10[49]);
AN2 GA10_50(oper2[50], oper1[10], g10[50]);
AN2 GA10_51(oper2[51], oper1[10], g10[51]);
AN2 GA10_52(oper2[52], oper1[10], g10[52]);
AN2 GA10_53(oper2[53], oper1[10], g10[53]);
AN2 GA10_54(oper2[54], oper1[10], g10[54]);
AN2 GA10_55(oper2[55], oper1[10], g10[55]);
AN2 GA10_56(oper2[56], oper1[10], g10[56]);
AN2 GA10_57(oper2[57], oper1[10], g10[57]);
AN2 GA10_58(oper2[58], oper1[10], g10[58]);
AN2 GA10_59(oper2[59], oper1[10], g10[59]);
AN2 GA10_60(oper2[60], oper1[10], g10[60]);
AN2 GA10_61(oper2[61], oper1[10], g10[61]);
AN2 GA10_62(oper2[62], oper1[10], g10[62]);
AN2 GA10_63(oper2[63], oper1[10], g10[63]);
AN2 GA9_8(oper2[8], oper1[9], g9[8]);
AN2 GA9_9(oper2[9], oper1[9], g9[9]);
AN2 GA9_10(oper2[10], oper1[9], g9[10]);
AN2 GA9_11(oper2[11], oper1[9], g9[11]);
AN2 GA9_12(oper2[12], oper1[9], g9[12]);
AN2 GA9_13(oper2[13], oper1[9], g9[13]);
AN2 GA9_14(oper2[14], oper1[9], g9[14]);
AN2 GA9_15(oper2[15], oper1[9], g9[15]);
AN2 GA9_16(oper2[16], oper1[9], g9[16]);
AN2 GA9_17(oper2[17], oper1[9], g9[17]);
AN2 GA9_18(oper2[18], oper1[9], g9[18]);
AN2 GA9_19(oper2[19], oper1[9], g9[19]);
AN2 GA9_20(oper2[20], oper1[9], g9[20]);
AN2 GA9_21(oper2[21], oper1[9], g9[21]);
AN2 GA9_22(oper2[22], oper1[9], g9[22]);
AN2 GA9_23(oper2[23], oper1[9], g9[23]);
AN2 GA9_24(oper2[24], oper1[9], g9[24]);
AN2 GA9_25(oper2[25], oper1[9], g9[25]);
AN2 GA9_26(oper2[26], oper1[9], g9[26]);
AN2 GA9_27(oper2[27], oper1[9], g9[27]);
AN2 GA9_28(oper2[28], oper1[9], g9[28]);
AN2 GA9_29(oper2[29], oper1[9], g9[29]);
AN2 GA9_30(oper2[30], oper1[9], g9[30]);
AN2 GA9_31(oper2[31], oper1[9], g9[31]);
AN2 GA9_32(oper2[32], oper1[9], g9[32]);
AN2 GA9_33(oper2[33], oper1[9], g9[33]);
AN2 GA9_34(oper2[34], oper1[9], g9[34]);
AN2 GA9_35(oper2[35], oper1[9], g9[35]);
AN2 GA9_36(oper2[36], oper1[9], g9[36]);
AN2 GA9_37(oper2[37], oper1[9], g9[37]);
AN2 GA9_38(oper2[38], oper1[9], g9[38]);
AN2 GA9_39(oper2[39], oper1[9], g9[39]);
AN2 GA9_40(oper2[40], oper1[9], g9[40]);
AN2 GA9_41(oper2[41], oper1[9], g9[41]);
AN2 GA9_42(oper2[42], oper1[9], g9[42]);
AN2 GA9_43(oper2[43], oper1[9], g9[43]);
AN2 GA9_44(oper2[44], oper1[9], g9[44]);
AN2 GA9_45(oper2[45], oper1[9], g9[45]);
AN2 GA9_46(oper2[46], oper1[9], g9[46]);
AN2 GA9_47(oper2[47], oper1[9], g9[47]);
AN2 GA9_48(oper2[48], oper1[9], g9[48]);
AN2 GA9_49(oper2[49], oper1[9], g9[49]);
AN2 GA9_50(oper2[50], oper1[9], g9[50]);
AN2 GA9_51(oper2[51], oper1[9], g9[51]);
AN2 GA9_52(oper2[52], oper1[9], g9[52]);
AN2 GA9_53(oper2[53], oper1[9], g9[53]);
AN2 GA9_54(oper2[54], oper1[9], g9[54]);
AN2 GA9_55(oper2[55], oper1[9], g9[55]);
AN2 GA9_56(oper2[56], oper1[9], g9[56]);
AN2 GA9_57(oper2[57], oper1[9], g9[57]);
AN2 GA9_58(oper2[58], oper1[9], g9[58]);
AN2 GA9_59(oper2[59], oper1[9], g9[59]);
AN2 GA9_60(oper2[60], oper1[9], g9[60]);
AN2 GA9_61(oper2[61], oper1[9], g9[61]);
AN2 GA9_62(oper2[62], oper1[9], g9[62]);
AN2 GA9_63(oper2[63], oper1[9], g9[63]);
AN2 GA8_8(oper2[8], oper1[8], g8[8]);
AN2 GA8_9(oper2[9], oper1[8], g8[9]);
AN2 GA8_10(oper2[10], oper1[8], g8[10]);
AN2 GA8_11(oper2[11], oper1[8], g8[11]);
AN2 GA8_12(oper2[12], oper1[8], g8[12]);
AN2 GA8_13(oper2[13], oper1[8], g8[13]);
AN2 GA8_14(oper2[14], oper1[8], g8[14]);
AN2 GA8_15(oper2[15], oper1[8], g8[15]);
AN2 GA8_16(oper2[16], oper1[8], g8[16]);
AN2 GA8_17(oper2[17], oper1[8], g8[17]);
AN2 GA8_18(oper2[18], oper1[8], g8[18]);
AN2 GA8_19(oper2[19], oper1[8], g8[19]);
AN2 GA8_20(oper2[20], oper1[8], g8[20]);
AN2 GA8_21(oper2[21], oper1[8], g8[21]);
AN2 GA8_22(oper2[22], oper1[8], g8[22]);
AN2 GA8_23(oper2[23], oper1[8], g8[23]);
AN2 GA8_24(oper2[24], oper1[8], g8[24]);
AN2 GA8_25(oper2[25], oper1[8], g8[25]);
AN2 GA8_26(oper2[26], oper1[8], g8[26]);
AN2 GA8_27(oper2[27], oper1[8], g8[27]);
AN2 GA8_28(oper2[28], oper1[8], g8[28]);
AN2 GA8_29(oper2[29], oper1[8], g8[29]);
AN2 GA8_30(oper2[30], oper1[8], g8[30]);
AN2 GA8_31(oper2[31], oper1[8], g8[31]);
AN2 GA8_32(oper2[32], oper1[8], g8[32]);
AN2 GA8_33(oper2[33], oper1[8], g8[33]);
AN2 GA8_34(oper2[34], oper1[8], g8[34]);
AN2 GA8_35(oper2[35], oper1[8], g8[35]);
AN2 GA8_36(oper2[36], oper1[8], g8[36]);
AN2 GA8_37(oper2[37], oper1[8], g8[37]);
AN2 GA8_38(oper2[38], oper1[8], g8[38]);
AN2 GA8_39(oper2[39], oper1[8], g8[39]);
AN2 GA8_40(oper2[40], oper1[8], g8[40]);
AN2 GA8_41(oper2[41], oper1[8], g8[41]);
AN2 GA8_42(oper2[42], oper1[8], g8[42]);
AN2 GA8_43(oper2[43], oper1[8], g8[43]);
AN2 GA8_44(oper2[44], oper1[8], g8[44]);
AN2 GA8_45(oper2[45], oper1[8], g8[45]);
AN2 GA8_46(oper2[46], oper1[8], g8[46]);
AN2 GA8_47(oper2[47], oper1[8], g8[47]);
AN2 GA8_48(oper2[48], oper1[8], g8[48]);
AN2 GA8_49(oper2[49], oper1[8], g8[49]);
AN2 GA8_50(oper2[50], oper1[8], g8[50]);
AN2 GA8_51(oper2[51], oper1[8], g8[51]);
AN2 GA8_52(oper2[52], oper1[8], g8[52]);
AN2 GA8_53(oper2[53], oper1[8], g8[53]);
AN2 GA8_54(oper2[54], oper1[8], g8[54]);
AN2 GA8_55(oper2[55], oper1[8], g8[55]);
AN2 GA8_56(oper2[56], oper1[8], g8[56]);
AN2 GA8_57(oper2[57], oper1[8], g8[57]);
AN2 GA8_58(oper2[58], oper1[8], g8[58]);
AN2 GA8_59(oper2[59], oper1[8], g8[59]);
AN2 GA8_60(oper2[60], oper1[8], g8[60]);
AN2 GA8_61(oper2[61], oper1[8], g8[61]);
AN2 GA8_62(oper2[62], oper1[8], g8[62]);
AN2 GA8_63(oper2[63], oper1[8], g8[63]);
FA1A GS62_9(g63[8], `zero, g62[9], ps62[9], pc62[9]);
FA1A GS62_10(g63[9], `zero, g62[10], ps62[10], pc62[10]);
FA1A GS62_11(g63[10], `zero, g62[11], ps62[11], pc62[11]);
FA1A GS62_12(g63[11], `zero, g62[12], ps62[12], pc62[12]);
FA1A GS62_13(g63[12], `zero, g62[13], ps62[13], pc62[13]);
FA1A GS62_14(g63[13], `zero, g62[14], ps62[14], pc62[14]);
FA1A GS62_15(g63[14], `zero, g62[15], ps62[15], pc62[15]);
FA1A GS62_16(g63[15], `zero, g62[16], ps62[16], pc62[16]);
FA1A GS62_17(g63[16], `zero, g62[17], ps62[17], pc62[17]);
FA1A GS62_18(g63[17], `zero, g62[18], ps62[18], pc62[18]);
FA1A GS62_19(g63[18], `zero, g62[19], ps62[19], pc62[19]);
FA1A GS62_20(g63[19], `zero, g62[20], ps62[20], pc62[20]);
FA1A GS62_21(g63[20], `zero, g62[21], ps62[21], pc62[21]);
FA1A GS62_22(g63[21], `zero, g62[22], ps62[22], pc62[22]);
FA1A GS62_23(g63[22], `zero, g62[23], ps62[23], pc62[23]);
FA1A GS62_24(g63[23], `zero, g62[24], ps62[24], pc62[24]);
FA1A GS62_25(g63[24], `zero, g62[25], ps62[25], pc62[25]);
FA1A GS62_26(g63[25], `zero, g62[26], ps62[26], pc62[26]);
FA1A GS62_27(g63[26], `zero, g62[27], ps62[27], pc62[27]);
FA1A GS62_28(g63[27], `zero, g62[28], ps62[28], pc62[28]);
FA1A GS62_29(g63[28], `zero, g62[29], ps62[29], pc62[29]);
FA1A GS62_30(g63[29], `zero, g62[30], ps62[30], pc62[30]);
FA1A GS62_31(g63[30], `zero, g62[31], ps62[31], pc62[31]);
FA1A GS62_32(g63[31], `zero, g62[32], ps62[32], pc62[32]);
FA1A GS62_33(g63[32], `zero, g62[33], ps62[33], pc62[33]);
FA1A GS62_34(g63[33], `zero, g62[34], ps62[34], pc62[34]);
FA1A GS62_35(g63[34], `zero, g62[35], ps62[35], pc62[35]);
FA1A GS62_36(g63[35], `zero, g62[36], ps62[36], pc62[36]);
FA1A GS62_37(g63[36], `zero, g62[37], ps62[37], pc62[37]);
FA1A GS62_38(g63[37], `zero, g62[38], ps62[38], pc62[38]);
FA1A GS62_39(g63[38], `zero, g62[39], ps62[39], pc62[39]);
FA1A GS62_40(g63[39], `zero, g62[40], ps62[40], pc62[40]);
FA1A GS62_41(g63[40], `zero, g62[41], ps62[41], pc62[41]);
FA1A GS62_42(g63[41], `zero, g62[42], ps62[42], pc62[42]);
FA1A GS62_43(g63[42], `zero, g62[43], ps62[43], pc62[43]);
FA1A GS62_44(g63[43], `zero, g62[44], ps62[44], pc62[44]);
FA1A GS62_45(g63[44], `zero, g62[45], ps62[45], pc62[45]);
FA1A GS62_46(g63[45], `zero, g62[46], ps62[46], pc62[46]);
FA1A GS62_47(g63[46], `zero, g62[47], ps62[47], pc62[47]);
FA1A GS62_48(g63[47], `zero, g62[48], ps62[48], pc62[48]);
FA1A GS62_49(g63[48], `zero, g62[49], ps62[49], pc62[49]);
FA1A GS62_50(g63[49], `zero, g62[50], ps62[50], pc62[50]);
FA1A GS62_51(g63[50], `zero, g62[51], ps62[51], pc62[51]);
FA1A GS62_52(g63[51], `zero, g62[52], ps62[52], pc62[52]);
FA1A GS62_53(g63[52], `zero, g62[53], ps62[53], pc62[53]);
FA1A GS62_54(g63[53], `zero, g62[54], ps62[54], pc62[54]);
FA1A GS62_55(g63[54], `zero, g62[55], ps62[55], pc62[55]);
FA1A GS62_56(g63[55], `zero, g62[56], ps62[56], pc62[56]);
FA1A GS62_57(g63[56], `zero, g62[57], ps62[57], pc62[57]);
FA1A GS62_58(g63[57], `zero, g62[58], ps62[58], pc62[58]);
FA1A GS62_59(g63[58], `zero, g62[59], ps62[59], pc62[59]);
FA1A GS62_60(g63[59], `zero, g62[60], ps62[60], pc62[60]);
FA1A GS62_61(g63[60], `zero, g62[61], ps62[61], pc62[61]);
FA1A GS62_62(g63[61], `zero, g62[62], ps62[62], pc62[62]);
FA1A GS62_63(g63[62], `zero, g62[63], ps62[63], pc62[63]);
FA1A GS61_9(g62[8], pc62[9], g61[9], ps61[9], pc61[9]);
FA1A GS61_10(ps62[9], pc62[10], g61[10], ps61[10], pc61[10]);
FA1A GS61_11(ps62[10], pc62[11], g61[11], ps61[11], pc61[11]);
FA1A GS61_12(ps62[11], pc62[12], g61[12], ps61[12], pc61[12]);
FA1A GS61_13(ps62[12], pc62[13], g61[13], ps61[13], pc61[13]);
FA1A GS61_14(ps62[13], pc62[14], g61[14], ps61[14], pc61[14]);
FA1A GS61_15(ps62[14], pc62[15], g61[15], ps61[15], pc61[15]);
FA1A GS61_16(ps62[15], pc62[16], g61[16], ps61[16], pc61[16]);
FA1A GS61_17(ps62[16], pc62[17], g61[17], ps61[17], pc61[17]);
FA1A GS61_18(ps62[17], pc62[18], g61[18], ps61[18], pc61[18]);
FA1A GS61_19(ps62[18], pc62[19], g61[19], ps61[19], pc61[19]);
FA1A GS61_20(ps62[19], pc62[20], g61[20], ps61[20], pc61[20]);
FA1A GS61_21(ps62[20], pc62[21], g61[21], ps61[21], pc61[21]);
FA1A GS61_22(ps62[21], pc62[22], g61[22], ps61[22], pc61[22]);
FA1A GS61_23(ps62[22], pc62[23], g61[23], ps61[23], pc61[23]);
FA1A GS61_24(ps62[23], pc62[24], g61[24], ps61[24], pc61[24]);
FA1A GS61_25(ps62[24], pc62[25], g61[25], ps61[25], pc61[25]);
FA1A GS61_26(ps62[25], pc62[26], g61[26], ps61[26], pc61[26]);
FA1A GS61_27(ps62[26], pc62[27], g61[27], ps61[27], pc61[27]);
FA1A GS61_28(ps62[27], pc62[28], g61[28], ps61[28], pc61[28]);
FA1A GS61_29(ps62[28], pc62[29], g61[29], ps61[29], pc61[29]);
FA1A GS61_30(ps62[29], pc62[30], g61[30], ps61[30], pc61[30]);
FA1A GS61_31(ps62[30], pc62[31], g61[31], ps61[31], pc61[31]);
FA1A GS61_32(ps62[31], pc62[32], g61[32], ps61[32], pc61[32]);
FA1A GS61_33(ps62[32], pc62[33], g61[33], ps61[33], pc61[33]);
FA1A GS61_34(ps62[33], pc62[34], g61[34], ps61[34], pc61[34]);
FA1A GS61_35(ps62[34], pc62[35], g61[35], ps61[35], pc61[35]);
FA1A GS61_36(ps62[35], pc62[36], g61[36], ps61[36], pc61[36]);
FA1A GS61_37(ps62[36], pc62[37], g61[37], ps61[37], pc61[37]);
FA1A GS61_38(ps62[37], pc62[38], g61[38], ps61[38], pc61[38]);
FA1A GS61_39(ps62[38], pc62[39], g61[39], ps61[39], pc61[39]);
FA1A GS61_40(ps62[39], pc62[40], g61[40], ps61[40], pc61[40]);
FA1A GS61_41(ps62[40], pc62[41], g61[41], ps61[41], pc61[41]);
FA1A GS61_42(ps62[41], pc62[42], g61[42], ps61[42], pc61[42]);
FA1A GS61_43(ps62[42], pc62[43], g61[43], ps61[43], pc61[43]);
FA1A GS61_44(ps62[43], pc62[44], g61[44], ps61[44], pc61[44]);
FA1A GS61_45(ps62[44], pc62[45], g61[45], ps61[45], pc61[45]);
FA1A GS61_46(ps62[45], pc62[46], g61[46], ps61[46], pc61[46]);
FA1A GS61_47(ps62[46], pc62[47], g61[47], ps61[47], pc61[47]);
FA1A GS61_48(ps62[47], pc62[48], g61[48], ps61[48], pc61[48]);
FA1A GS61_49(ps62[48], pc62[49], g61[49], ps61[49], pc61[49]);
FA1A GS61_50(ps62[49], pc62[50], g61[50], ps61[50], pc61[50]);
FA1A GS61_51(ps62[50], pc62[51], g61[51], ps61[51], pc61[51]);
FA1A GS61_52(ps62[51], pc62[52], g61[52], ps61[52], pc61[52]);
FA1A GS61_53(ps62[52], pc62[53], g61[53], ps61[53], pc61[53]);
FA1A GS61_54(ps62[53], pc62[54], g61[54], ps61[54], pc61[54]);
FA1A GS61_55(ps62[54], pc62[55], g61[55], ps61[55], pc61[55]);
FA1A GS61_56(ps62[55], pc62[56], g61[56], ps61[56], pc61[56]);
FA1A GS61_57(ps62[56], pc62[57], g61[57], ps61[57], pc61[57]);
FA1A GS61_58(ps62[57], pc62[58], g61[58], ps61[58], pc61[58]);
FA1A GS61_59(ps62[58], pc62[59], g61[59], ps61[59], pc61[59]);
FA1A GS61_60(ps62[59], pc62[60], g61[60], ps61[60], pc61[60]);
FA1A GS61_61(ps62[60], pc62[61], g61[61], ps61[61], pc61[61]);
FA1A GS61_62(ps62[61], pc62[62], g61[62], ps61[62], pc61[62]);
FA1A GS61_63(ps62[62], pc62[63], g61[63], ps61[63], pc61[63]);
FA1A GS60_9(g61[8], pc61[9], g60[9], ps60[9], pc60[9]);
FA1A GS60_10(ps61[9], pc61[10], g60[10], ps60[10], pc60[10]);
FA1A GS60_11(ps61[10], pc61[11], g60[11], ps60[11], pc60[11]);
FA1A GS60_12(ps61[11], pc61[12], g60[12], ps60[12], pc60[12]);
FA1A GS60_13(ps61[12], pc61[13], g60[13], ps60[13], pc60[13]);
FA1A GS60_14(ps61[13], pc61[14], g60[14], ps60[14], pc60[14]);
FA1A GS60_15(ps61[14], pc61[15], g60[15], ps60[15], pc60[15]);
FA1A GS60_16(ps61[15], pc61[16], g60[16], ps60[16], pc60[16]);
FA1A GS60_17(ps61[16], pc61[17], g60[17], ps60[17], pc60[17]);
FA1A GS60_18(ps61[17], pc61[18], g60[18], ps60[18], pc60[18]);
FA1A GS60_19(ps61[18], pc61[19], g60[19], ps60[19], pc60[19]);
FA1A GS60_20(ps61[19], pc61[20], g60[20], ps60[20], pc60[20]);
FA1A GS60_21(ps61[20], pc61[21], g60[21], ps60[21], pc60[21]);
FA1A GS60_22(ps61[21], pc61[22], g60[22], ps60[22], pc60[22]);
FA1A GS60_23(ps61[22], pc61[23], g60[23], ps60[23], pc60[23]);
FA1A GS60_24(ps61[23], pc61[24], g60[24], ps60[24], pc60[24]);
FA1A GS60_25(ps61[24], pc61[25], g60[25], ps60[25], pc60[25]);
FA1A GS60_26(ps61[25], pc61[26], g60[26], ps60[26], pc60[26]);
FA1A GS60_27(ps61[26], pc61[27], g60[27], ps60[27], pc60[27]);
FA1A GS60_28(ps61[27], pc61[28], g60[28], ps60[28], pc60[28]);
FA1A GS60_29(ps61[28], pc61[29], g60[29], ps60[29], pc60[29]);
FA1A GS60_30(ps61[29], pc61[30], g60[30], ps60[30], pc60[30]);
FA1A GS60_31(ps61[30], pc61[31], g60[31], ps60[31], pc60[31]);
FA1A GS60_32(ps61[31], pc61[32], g60[32], ps60[32], pc60[32]);
FA1A GS60_33(ps61[32], pc61[33], g60[33], ps60[33], pc60[33]);
FA1A GS60_34(ps61[33], pc61[34], g60[34], ps60[34], pc60[34]);
FA1A GS60_35(ps61[34], pc61[35], g60[35], ps60[35], pc60[35]);
FA1A GS60_36(ps61[35], pc61[36], g60[36], ps60[36], pc60[36]);
FA1A GS60_37(ps61[36], pc61[37], g60[37], ps60[37], pc60[37]);
FA1A GS60_38(ps61[37], pc61[38], g60[38], ps60[38], pc60[38]);
FA1A GS60_39(ps61[38], pc61[39], g60[39], ps60[39], pc60[39]);
FA1A GS60_40(ps61[39], pc61[40], g60[40], ps60[40], pc60[40]);
FA1A GS60_41(ps61[40], pc61[41], g60[41], ps60[41], pc60[41]);
FA1A GS60_42(ps61[41], pc61[42], g60[42], ps60[42], pc60[42]);
FA1A GS60_43(ps61[42], pc61[43], g60[43], ps60[43], pc60[43]);
FA1A GS60_44(ps61[43], pc61[44], g60[44], ps60[44], pc60[44]);
FA1A GS60_45(ps61[44], pc61[45], g60[45], ps60[45], pc60[45]);
FA1A GS60_46(ps61[45], pc61[46], g60[46], ps60[46], pc60[46]);
FA1A GS60_47(ps61[46], pc61[47], g60[47], ps60[47], pc60[47]);
FA1A GS60_48(ps61[47], pc61[48], g60[48], ps60[48], pc60[48]);
FA1A GS60_49(ps61[48], pc61[49], g60[49], ps60[49], pc60[49]);
FA1A GS60_50(ps61[49], pc61[50], g60[50], ps60[50], pc60[50]);
FA1A GS60_51(ps61[50], pc61[51], g60[51], ps60[51], pc60[51]);
FA1A GS60_52(ps61[51], pc61[52], g60[52], ps60[52], pc60[52]);
FA1A GS60_53(ps61[52], pc61[53], g60[53], ps60[53], pc60[53]);
FA1A GS60_54(ps61[53], pc61[54], g60[54], ps60[54], pc60[54]);
FA1A GS60_55(ps61[54], pc61[55], g60[55], ps60[55], pc60[55]);
FA1A GS60_56(ps61[55], pc61[56], g60[56], ps60[56], pc60[56]);
FA1A GS60_57(ps61[56], pc61[57], g60[57], ps60[57], pc60[57]);
FA1A GS60_58(ps61[57], pc61[58], g60[58], ps60[58], pc60[58]);
FA1A GS60_59(ps61[58], pc61[59], g60[59], ps60[59], pc60[59]);
FA1A GS60_60(ps61[59], pc61[60], g60[60], ps60[60], pc60[60]);
FA1A GS60_61(ps61[60], pc61[61], g60[61], ps60[61], pc60[61]);
FA1A GS60_62(ps61[61], pc61[62], g60[62], ps60[62], pc60[62]);
FA1A GS60_63(ps61[62], pc61[63], g60[63], ps60[63], pc60[63]);
FA1A GS59_9(g60[8], pc60[9], g59[9], ps59[9], pc59[9]);
FA1A GS59_10(ps60[9], pc60[10], g59[10], ps59[10], pc59[10]);
FA1A GS59_11(ps60[10], pc60[11], g59[11], ps59[11], pc59[11]);
FA1A GS59_12(ps60[11], pc60[12], g59[12], ps59[12], pc59[12]);
FA1A GS59_13(ps60[12], pc60[13], g59[13], ps59[13], pc59[13]);
FA1A GS59_14(ps60[13], pc60[14], g59[14], ps59[14], pc59[14]);
FA1A GS59_15(ps60[14], pc60[15], g59[15], ps59[15], pc59[15]);
FA1A GS59_16(ps60[15], pc60[16], g59[16], ps59[16], pc59[16]);
FA1A GS59_17(ps60[16], pc60[17], g59[17], ps59[17], pc59[17]);
FA1A GS59_18(ps60[17], pc60[18], g59[18], ps59[18], pc59[18]);
FA1A GS59_19(ps60[18], pc60[19], g59[19], ps59[19], pc59[19]);
FA1A GS59_20(ps60[19], pc60[20], g59[20], ps59[20], pc59[20]);
FA1A GS59_21(ps60[20], pc60[21], g59[21], ps59[21], pc59[21]);
FA1A GS59_22(ps60[21], pc60[22], g59[22], ps59[22], pc59[22]);
FA1A GS59_23(ps60[22], pc60[23], g59[23], ps59[23], pc59[23]);
FA1A GS59_24(ps60[23], pc60[24], g59[24], ps59[24], pc59[24]);
FA1A GS59_25(ps60[24], pc60[25], g59[25], ps59[25], pc59[25]);
FA1A GS59_26(ps60[25], pc60[26], g59[26], ps59[26], pc59[26]);
FA1A GS59_27(ps60[26], pc60[27], g59[27], ps59[27], pc59[27]);
FA1A GS59_28(ps60[27], pc60[28], g59[28], ps59[28], pc59[28]);
FA1A GS59_29(ps60[28], pc60[29], g59[29], ps59[29], pc59[29]);
FA1A GS59_30(ps60[29], pc60[30], g59[30], ps59[30], pc59[30]);
FA1A GS59_31(ps60[30], pc60[31], g59[31], ps59[31], pc59[31]);
FA1A GS59_32(ps60[31], pc60[32], g59[32], ps59[32], pc59[32]);
FA1A GS59_33(ps60[32], pc60[33], g59[33], ps59[33], pc59[33]);
FA1A GS59_34(ps60[33], pc60[34], g59[34], ps59[34], pc59[34]);
FA1A GS59_35(ps60[34], pc60[35], g59[35], ps59[35], pc59[35]);
FA1A GS59_36(ps60[35], pc60[36], g59[36], ps59[36], pc59[36]);
FA1A GS59_37(ps60[36], pc60[37], g59[37], ps59[37], pc59[37]);
FA1A GS59_38(ps60[37], pc60[38], g59[38], ps59[38], pc59[38]);
FA1A GS59_39(ps60[38], pc60[39], g59[39], ps59[39], pc59[39]);
FA1A GS59_40(ps60[39], pc60[40], g59[40], ps59[40], pc59[40]);
FA1A GS59_41(ps60[40], pc60[41], g59[41], ps59[41], pc59[41]);
FA1A GS59_42(ps60[41], pc60[42], g59[42], ps59[42], pc59[42]);
FA1A GS59_43(ps60[42], pc60[43], g59[43], ps59[43], pc59[43]);
FA1A GS59_44(ps60[43], pc60[44], g59[44], ps59[44], pc59[44]);
FA1A GS59_45(ps60[44], pc60[45], g59[45], ps59[45], pc59[45]);
FA1A GS59_46(ps60[45], pc60[46], g59[46], ps59[46], pc59[46]);
FA1A GS59_47(ps60[46], pc60[47], g59[47], ps59[47], pc59[47]);
FA1A GS59_48(ps60[47], pc60[48], g59[48], ps59[48], pc59[48]);
FA1A GS59_49(ps60[48], pc60[49], g59[49], ps59[49], pc59[49]);
FA1A GS59_50(ps60[49], pc60[50], g59[50], ps59[50], pc59[50]);
FA1A GS59_51(ps60[50], pc60[51], g59[51], ps59[51], pc59[51]);
FA1A GS59_52(ps60[51], pc60[52], g59[52], ps59[52], pc59[52]);
FA1A GS59_53(ps60[52], pc60[53], g59[53], ps59[53], pc59[53]);
FA1A GS59_54(ps60[53], pc60[54], g59[54], ps59[54], pc59[54]);
FA1A GS59_55(ps60[54], pc60[55], g59[55], ps59[55], pc59[55]);
FA1A GS59_56(ps60[55], pc60[56], g59[56], ps59[56], pc59[56]);
FA1A GS59_57(ps60[56], pc60[57], g59[57], ps59[57], pc59[57]);
FA1A GS59_58(ps60[57], pc60[58], g59[58], ps59[58], pc59[58]);
FA1A GS59_59(ps60[58], pc60[59], g59[59], ps59[59], pc59[59]);
FA1A GS59_60(ps60[59], pc60[60], g59[60], ps59[60], pc59[60]);
FA1A GS59_61(ps60[60], pc60[61], g59[61], ps59[61], pc59[61]);
FA1A GS59_62(ps60[61], pc60[62], g59[62], ps59[62], pc59[62]);
FA1A GS59_63(ps60[62], pc60[63], g59[63], ps59[63], pc59[63]);
FA1A GS58_9(g59[8], pc59[9], g58[9], ps58[9], pc58[9]);
FA1A GS58_10(ps59[9], pc59[10], g58[10], ps58[10], pc58[10]);
FA1A GS58_11(ps59[10], pc59[11], g58[11], ps58[11], pc58[11]);
FA1A GS58_12(ps59[11], pc59[12], g58[12], ps58[12], pc58[12]);
FA1A GS58_13(ps59[12], pc59[13], g58[13], ps58[13], pc58[13]);
FA1A GS58_14(ps59[13], pc59[14], g58[14], ps58[14], pc58[14]);
FA1A GS58_15(ps59[14], pc59[15], g58[15], ps58[15], pc58[15]);
FA1A GS58_16(ps59[15], pc59[16], g58[16], ps58[16], pc58[16]);
FA1A GS58_17(ps59[16], pc59[17], g58[17], ps58[17], pc58[17]);
FA1A GS58_18(ps59[17], pc59[18], g58[18], ps58[18], pc58[18]);
FA1A GS58_19(ps59[18], pc59[19], g58[19], ps58[19], pc58[19]);
FA1A GS58_20(ps59[19], pc59[20], g58[20], ps58[20], pc58[20]);
FA1A GS58_21(ps59[20], pc59[21], g58[21], ps58[21], pc58[21]);
FA1A GS58_22(ps59[21], pc59[22], g58[22], ps58[22], pc58[22]);
FA1A GS58_23(ps59[22], pc59[23], g58[23], ps58[23], pc58[23]);
FA1A GS58_24(ps59[23], pc59[24], g58[24], ps58[24], pc58[24]);
FA1A GS58_25(ps59[24], pc59[25], g58[25], ps58[25], pc58[25]);
FA1A GS58_26(ps59[25], pc59[26], g58[26], ps58[26], pc58[26]);
FA1A GS58_27(ps59[26], pc59[27], g58[27], ps58[27], pc58[27]);
FA1A GS58_28(ps59[27], pc59[28], g58[28], ps58[28], pc58[28]);
FA1A GS58_29(ps59[28], pc59[29], g58[29], ps58[29], pc58[29]);
FA1A GS58_30(ps59[29], pc59[30], g58[30], ps58[30], pc58[30]);
FA1A GS58_31(ps59[30], pc59[31], g58[31], ps58[31], pc58[31]);
FA1A GS58_32(ps59[31], pc59[32], g58[32], ps58[32], pc58[32]);
FA1A GS58_33(ps59[32], pc59[33], g58[33], ps58[33], pc58[33]);
FA1A GS58_34(ps59[33], pc59[34], g58[34], ps58[34], pc58[34]);
FA1A GS58_35(ps59[34], pc59[35], g58[35], ps58[35], pc58[35]);
FA1A GS58_36(ps59[35], pc59[36], g58[36], ps58[36], pc58[36]);
FA1A GS58_37(ps59[36], pc59[37], g58[37], ps58[37], pc58[37]);
FA1A GS58_38(ps59[37], pc59[38], g58[38], ps58[38], pc58[38]);
FA1A GS58_39(ps59[38], pc59[39], g58[39], ps58[39], pc58[39]);
FA1A GS58_40(ps59[39], pc59[40], g58[40], ps58[40], pc58[40]);
FA1A GS58_41(ps59[40], pc59[41], g58[41], ps58[41], pc58[41]);
FA1A GS58_42(ps59[41], pc59[42], g58[42], ps58[42], pc58[42]);
FA1A GS58_43(ps59[42], pc59[43], g58[43], ps58[43], pc58[43]);
FA1A GS58_44(ps59[43], pc59[44], g58[44], ps58[44], pc58[44]);
FA1A GS58_45(ps59[44], pc59[45], g58[45], ps58[45], pc58[45]);
FA1A GS58_46(ps59[45], pc59[46], g58[46], ps58[46], pc58[46]);
FA1A GS58_47(ps59[46], pc59[47], g58[47], ps58[47], pc58[47]);
FA1A GS58_48(ps59[47], pc59[48], g58[48], ps58[48], pc58[48]);
FA1A GS58_49(ps59[48], pc59[49], g58[49], ps58[49], pc58[49]);
FA1A GS58_50(ps59[49], pc59[50], g58[50], ps58[50], pc58[50]);
FA1A GS58_51(ps59[50], pc59[51], g58[51], ps58[51], pc58[51]);
FA1A GS58_52(ps59[51], pc59[52], g58[52], ps58[52], pc58[52]);
FA1A GS58_53(ps59[52], pc59[53], g58[53], ps58[53], pc58[53]);
FA1A GS58_54(ps59[53], pc59[54], g58[54], ps58[54], pc58[54]);
FA1A GS58_55(ps59[54], pc59[55], g58[55], ps58[55], pc58[55]);
FA1A GS58_56(ps59[55], pc59[56], g58[56], ps58[56], pc58[56]);
FA1A GS58_57(ps59[56], pc59[57], g58[57], ps58[57], pc58[57]);
FA1A GS58_58(ps59[57], pc59[58], g58[58], ps58[58], pc58[58]);
FA1A GS58_59(ps59[58], pc59[59], g58[59], ps58[59], pc58[59]);
FA1A GS58_60(ps59[59], pc59[60], g58[60], ps58[60], pc58[60]);
FA1A GS58_61(ps59[60], pc59[61], g58[61], ps58[61], pc58[61]);
FA1A GS58_62(ps59[61], pc59[62], g58[62], ps58[62], pc58[62]);
FA1A GS58_63(ps59[62], pc59[63], g58[63], ps58[63], pc58[63]);
FA1A GS57_9(g58[8], pc58[9], g57[9], ps57[9], pc57[9]);
FA1A GS57_10(ps58[9], pc58[10], g57[10], ps57[10], pc57[10]);
FA1A GS57_11(ps58[10], pc58[11], g57[11], ps57[11], pc57[11]);
FA1A GS57_12(ps58[11], pc58[12], g57[12], ps57[12], pc57[12]);
FA1A GS57_13(ps58[12], pc58[13], g57[13], ps57[13], pc57[13]);
FA1A GS57_14(ps58[13], pc58[14], g57[14], ps57[14], pc57[14]);
FA1A GS57_15(ps58[14], pc58[15], g57[15], ps57[15], pc57[15]);
FA1A GS57_16(ps58[15], pc58[16], g57[16], ps57[16], pc57[16]);
FA1A GS57_17(ps58[16], pc58[17], g57[17], ps57[17], pc57[17]);
FA1A GS57_18(ps58[17], pc58[18], g57[18], ps57[18], pc57[18]);
FA1A GS57_19(ps58[18], pc58[19], g57[19], ps57[19], pc57[19]);
FA1A GS57_20(ps58[19], pc58[20], g57[20], ps57[20], pc57[20]);
FA1A GS57_21(ps58[20], pc58[21], g57[21], ps57[21], pc57[21]);
FA1A GS57_22(ps58[21], pc58[22], g57[22], ps57[22], pc57[22]);
FA1A GS57_23(ps58[22], pc58[23], g57[23], ps57[23], pc57[23]);
FA1A GS57_24(ps58[23], pc58[24], g57[24], ps57[24], pc57[24]);
FA1A GS57_25(ps58[24], pc58[25], g57[25], ps57[25], pc57[25]);
FA1A GS57_26(ps58[25], pc58[26], g57[26], ps57[26], pc57[26]);
FA1A GS57_27(ps58[26], pc58[27], g57[27], ps57[27], pc57[27]);
FA1A GS57_28(ps58[27], pc58[28], g57[28], ps57[28], pc57[28]);
FA1A GS57_29(ps58[28], pc58[29], g57[29], ps57[29], pc57[29]);
FA1A GS57_30(ps58[29], pc58[30], g57[30], ps57[30], pc57[30]);
FA1A GS57_31(ps58[30], pc58[31], g57[31], ps57[31], pc57[31]);
FA1A GS57_32(ps58[31], pc58[32], g57[32], ps57[32], pc57[32]);
FA1A GS57_33(ps58[32], pc58[33], g57[33], ps57[33], pc57[33]);
FA1A GS57_34(ps58[33], pc58[34], g57[34], ps57[34], pc57[34]);
FA1A GS57_35(ps58[34], pc58[35], g57[35], ps57[35], pc57[35]);
FA1A GS57_36(ps58[35], pc58[36], g57[36], ps57[36], pc57[36]);
FA1A GS57_37(ps58[36], pc58[37], g57[37], ps57[37], pc57[37]);
FA1A GS57_38(ps58[37], pc58[38], g57[38], ps57[38], pc57[38]);
FA1A GS57_39(ps58[38], pc58[39], g57[39], ps57[39], pc57[39]);
FA1A GS57_40(ps58[39], pc58[40], g57[40], ps57[40], pc57[40]);
FA1A GS57_41(ps58[40], pc58[41], g57[41], ps57[41], pc57[41]);
FA1A GS57_42(ps58[41], pc58[42], g57[42], ps57[42], pc57[42]);
FA1A GS57_43(ps58[42], pc58[43], g57[43], ps57[43], pc57[43]);
FA1A GS57_44(ps58[43], pc58[44], g57[44], ps57[44], pc57[44]);
FA1A GS57_45(ps58[44], pc58[45], g57[45], ps57[45], pc57[45]);
FA1A GS57_46(ps58[45], pc58[46], g57[46], ps57[46], pc57[46]);
FA1A GS57_47(ps58[46], pc58[47], g57[47], ps57[47], pc57[47]);
FA1A GS57_48(ps58[47], pc58[48], g57[48], ps57[48], pc57[48]);
FA1A GS57_49(ps58[48], pc58[49], g57[49], ps57[49], pc57[49]);
FA1A GS57_50(ps58[49], pc58[50], g57[50], ps57[50], pc57[50]);
FA1A GS57_51(ps58[50], pc58[51], g57[51], ps57[51], pc57[51]);
FA1A GS57_52(ps58[51], pc58[52], g57[52], ps57[52], pc57[52]);
FA1A GS57_53(ps58[52], pc58[53], g57[53], ps57[53], pc57[53]);
FA1A GS57_54(ps58[53], pc58[54], g57[54], ps57[54], pc57[54]);
FA1A GS57_55(ps58[54], pc58[55], g57[55], ps57[55], pc57[55]);
FA1A GS57_56(ps58[55], pc58[56], g57[56], ps57[56], pc57[56]);
FA1A GS57_57(ps58[56], pc58[57], g57[57], ps57[57], pc57[57]);
FA1A GS57_58(ps58[57], pc58[58], g57[58], ps57[58], pc57[58]);
FA1A GS57_59(ps58[58], pc58[59], g57[59], ps57[59], pc57[59]);
FA1A GS57_60(ps58[59], pc58[60], g57[60], ps57[60], pc57[60]);
FA1A GS57_61(ps58[60], pc58[61], g57[61], ps57[61], pc57[61]);
FA1A GS57_62(ps58[61], pc58[62], g57[62], ps57[62], pc57[62]);
FA1A GS57_63(ps58[62], pc58[63], g57[63], ps57[63], pc57[63]);
FA1A GS56_9(g57[8], pc57[9], g56[9], ps56[9], pc56[9]);
FA1A GS56_10(ps57[9], pc57[10], g56[10], ps56[10], pc56[10]);
FA1A GS56_11(ps57[10], pc57[11], g56[11], ps56[11], pc56[11]);
FA1A GS56_12(ps57[11], pc57[12], g56[12], ps56[12], pc56[12]);
FA1A GS56_13(ps57[12], pc57[13], g56[13], ps56[13], pc56[13]);
FA1A GS56_14(ps57[13], pc57[14], g56[14], ps56[14], pc56[14]);
FA1A GS56_15(ps57[14], pc57[15], g56[15], ps56[15], pc56[15]);
FA1A GS56_16(ps57[15], pc57[16], g56[16], ps56[16], pc56[16]);
FA1A GS56_17(ps57[16], pc57[17], g56[17], ps56[17], pc56[17]);
FA1A GS56_18(ps57[17], pc57[18], g56[18], ps56[18], pc56[18]);
FA1A GS56_19(ps57[18], pc57[19], g56[19], ps56[19], pc56[19]);
FA1A GS56_20(ps57[19], pc57[20], g56[20], ps56[20], pc56[20]);
FA1A GS56_21(ps57[20], pc57[21], g56[21], ps56[21], pc56[21]);
FA1A GS56_22(ps57[21], pc57[22], g56[22], ps56[22], pc56[22]);
FA1A GS56_23(ps57[22], pc57[23], g56[23], ps56[23], pc56[23]);
FA1A GS56_24(ps57[23], pc57[24], g56[24], ps56[24], pc56[24]);
FA1A GS56_25(ps57[24], pc57[25], g56[25], ps56[25], pc56[25]);
FA1A GS56_26(ps57[25], pc57[26], g56[26], ps56[26], pc56[26]);
FA1A GS56_27(ps57[26], pc57[27], g56[27], ps56[27], pc56[27]);
FA1A GS56_28(ps57[27], pc57[28], g56[28], ps56[28], pc56[28]);
FA1A GS56_29(ps57[28], pc57[29], g56[29], ps56[29], pc56[29]);
FA1A GS56_30(ps57[29], pc57[30], g56[30], ps56[30], pc56[30]);
FA1A GS56_31(ps57[30], pc57[31], g56[31], ps56[31], pc56[31]);
FA1A GS56_32(ps57[31], pc57[32], g56[32], ps56[32], pc56[32]);
FA1A GS56_33(ps57[32], pc57[33], g56[33], ps56[33], pc56[33]);
FA1A GS56_34(ps57[33], pc57[34], g56[34], ps56[34], pc56[34]);
FA1A GS56_35(ps57[34], pc57[35], g56[35], ps56[35], pc56[35]);
FA1A GS56_36(ps57[35], pc57[36], g56[36], ps56[36], pc56[36]);
FA1A GS56_37(ps57[36], pc57[37], g56[37], ps56[37], pc56[37]);
FA1A GS56_38(ps57[37], pc57[38], g56[38], ps56[38], pc56[38]);
FA1A GS56_39(ps57[38], pc57[39], g56[39], ps56[39], pc56[39]);
FA1A GS56_40(ps57[39], pc57[40], g56[40], ps56[40], pc56[40]);
FA1A GS56_41(ps57[40], pc57[41], g56[41], ps56[41], pc56[41]);
FA1A GS56_42(ps57[41], pc57[42], g56[42], ps56[42], pc56[42]);
FA1A GS56_43(ps57[42], pc57[43], g56[43], ps56[43], pc56[43]);
FA1A GS56_44(ps57[43], pc57[44], g56[44], ps56[44], pc56[44]);
FA1A GS56_45(ps57[44], pc57[45], g56[45], ps56[45], pc56[45]);
FA1A GS56_46(ps57[45], pc57[46], g56[46], ps56[46], pc56[46]);
FA1A GS56_47(ps57[46], pc57[47], g56[47], ps56[47], pc56[47]);
FA1A GS56_48(ps57[47], pc57[48], g56[48], ps56[48], pc56[48]);
FA1A GS56_49(ps57[48], pc57[49], g56[49], ps56[49], pc56[49]);
FA1A GS56_50(ps57[49], pc57[50], g56[50], ps56[50], pc56[50]);
FA1A GS56_51(ps57[50], pc57[51], g56[51], ps56[51], pc56[51]);
FA1A GS56_52(ps57[51], pc57[52], g56[52], ps56[52], pc56[52]);
FA1A GS56_53(ps57[52], pc57[53], g56[53], ps56[53], pc56[53]);
FA1A GS56_54(ps57[53], pc57[54], g56[54], ps56[54], pc56[54]);
FA1A GS56_55(ps57[54], pc57[55], g56[55], ps56[55], pc56[55]);
FA1A GS56_56(ps57[55], pc57[56], g56[56], ps56[56], pc56[56]);
FA1A GS56_57(ps57[56], pc57[57], g56[57], ps56[57], pc56[57]);
FA1A GS56_58(ps57[57], pc57[58], g56[58], ps56[58], pc56[58]);
FA1A GS56_59(ps57[58], pc57[59], g56[59], ps56[59], pc56[59]);
FA1A GS56_60(ps57[59], pc57[60], g56[60], ps56[60], pc56[60]);
FA1A GS56_61(ps57[60], pc57[61], g56[61], ps56[61], pc56[61]);
FA1A GS56_62(ps57[61], pc57[62], g56[62], ps56[62], pc56[62]);
FA1A GS56_63(ps57[62], pc57[63], g56[63], ps56[63], pc56[63]);
FA1A GS55_9(g56[8], pc56[9], g55[9], ps55[9], pc55[9]);
FA1A GS55_10(ps56[9], pc56[10], g55[10], ps55[10], pc55[10]);
FA1A GS55_11(ps56[10], pc56[11], g55[11], ps55[11], pc55[11]);
FA1A GS55_12(ps56[11], pc56[12], g55[12], ps55[12], pc55[12]);
FA1A GS55_13(ps56[12], pc56[13], g55[13], ps55[13], pc55[13]);
FA1A GS55_14(ps56[13], pc56[14], g55[14], ps55[14], pc55[14]);
FA1A GS55_15(ps56[14], pc56[15], g55[15], ps55[15], pc55[15]);
FA1A GS55_16(ps56[15], pc56[16], g55[16], ps55[16], pc55[16]);
FA1A GS55_17(ps56[16], pc56[17], g55[17], ps55[17], pc55[17]);
FA1A GS55_18(ps56[17], pc56[18], g55[18], ps55[18], pc55[18]);
FA1A GS55_19(ps56[18], pc56[19], g55[19], ps55[19], pc55[19]);
FA1A GS55_20(ps56[19], pc56[20], g55[20], ps55[20], pc55[20]);
FA1A GS55_21(ps56[20], pc56[21], g55[21], ps55[21], pc55[21]);
FA1A GS55_22(ps56[21], pc56[22], g55[22], ps55[22], pc55[22]);
FA1A GS55_23(ps56[22], pc56[23], g55[23], ps55[23], pc55[23]);
FA1A GS55_24(ps56[23], pc56[24], g55[24], ps55[24], pc55[24]);
FA1A GS55_25(ps56[24], pc56[25], g55[25], ps55[25], pc55[25]);
FA1A GS55_26(ps56[25], pc56[26], g55[26], ps55[26], pc55[26]);
FA1A GS55_27(ps56[26], pc56[27], g55[27], ps55[27], pc55[27]);
FA1A GS55_28(ps56[27], pc56[28], g55[28], ps55[28], pc55[28]);
FA1A GS55_29(ps56[28], pc56[29], g55[29], ps55[29], pc55[29]);
FA1A GS55_30(ps56[29], pc56[30], g55[30], ps55[30], pc55[30]);
FA1A GS55_31(ps56[30], pc56[31], g55[31], ps55[31], pc55[31]);
FA1A GS55_32(ps56[31], pc56[32], g55[32], ps55[32], pc55[32]);
FA1A GS55_33(ps56[32], pc56[33], g55[33], ps55[33], pc55[33]);
FA1A GS55_34(ps56[33], pc56[34], g55[34], ps55[34], pc55[34]);
FA1A GS55_35(ps56[34], pc56[35], g55[35], ps55[35], pc55[35]);
FA1A GS55_36(ps56[35], pc56[36], g55[36], ps55[36], pc55[36]);
FA1A GS55_37(ps56[36], pc56[37], g55[37], ps55[37], pc55[37]);
FA1A GS55_38(ps56[37], pc56[38], g55[38], ps55[38], pc55[38]);
FA1A GS55_39(ps56[38], pc56[39], g55[39], ps55[39], pc55[39]);
FA1A GS55_40(ps56[39], pc56[40], g55[40], ps55[40], pc55[40]);
FA1A GS55_41(ps56[40], pc56[41], g55[41], ps55[41], pc55[41]);
FA1A GS55_42(ps56[41], pc56[42], g55[42], ps55[42], pc55[42]);
FA1A GS55_43(ps56[42], pc56[43], g55[43], ps55[43], pc55[43]);
FA1A GS55_44(ps56[43], pc56[44], g55[44], ps55[44], pc55[44]);
FA1A GS55_45(ps56[44], pc56[45], g55[45], ps55[45], pc55[45]);
FA1A GS55_46(ps56[45], pc56[46], g55[46], ps55[46], pc55[46]);
FA1A GS55_47(ps56[46], pc56[47], g55[47], ps55[47], pc55[47]);
FA1A GS55_48(ps56[47], pc56[48], g55[48], ps55[48], pc55[48]);
FA1A GS55_49(ps56[48], pc56[49], g55[49], ps55[49], pc55[49]);
FA1A GS55_50(ps56[49], pc56[50], g55[50], ps55[50], pc55[50]);
FA1A GS55_51(ps56[50], pc56[51], g55[51], ps55[51], pc55[51]);
FA1A GS55_52(ps56[51], pc56[52], g55[52], ps55[52], pc55[52]);
FA1A GS55_53(ps56[52], pc56[53], g55[53], ps55[53], pc55[53]);
FA1A GS55_54(ps56[53], pc56[54], g55[54], ps55[54], pc55[54]);
FA1A GS55_55(ps56[54], pc56[55], g55[55], ps55[55], pc55[55]);
FA1A GS55_56(ps56[55], pc56[56], g55[56], ps55[56], pc55[56]);
FA1A GS55_57(ps56[56], pc56[57], g55[57], ps55[57], pc55[57]);
FA1A GS55_58(ps56[57], pc56[58], g55[58], ps55[58], pc55[58]);
FA1A GS55_59(ps56[58], pc56[59], g55[59], ps55[59], pc55[59]);
FA1A GS55_60(ps56[59], pc56[60], g55[60], ps55[60], pc55[60]);
FA1A GS55_61(ps56[60], pc56[61], g55[61], ps55[61], pc55[61]);
FA1A GS55_62(ps56[61], pc56[62], g55[62], ps55[62], pc55[62]);
FA1A GS55_63(ps56[62], pc56[63], g55[63], ps55[63], pc55[63]);
FA1A GS54_9(g55[8], pc55[9], g54[9], ps54[9], pc54[9]);
FA1A GS54_10(ps55[9], pc55[10], g54[10], ps54[10], pc54[10]);
FA1A GS54_11(ps55[10], pc55[11], g54[11], ps54[11], pc54[11]);
FA1A GS54_12(ps55[11], pc55[12], g54[12], ps54[12], pc54[12]);
FA1A GS54_13(ps55[12], pc55[13], g54[13], ps54[13], pc54[13]);
FA1A GS54_14(ps55[13], pc55[14], g54[14], ps54[14], pc54[14]);
FA1A GS54_15(ps55[14], pc55[15], g54[15], ps54[15], pc54[15]);
FA1A GS54_16(ps55[15], pc55[16], g54[16], ps54[16], pc54[16]);
FA1A GS54_17(ps55[16], pc55[17], g54[17], ps54[17], pc54[17]);
FA1A GS54_18(ps55[17], pc55[18], g54[18], ps54[18], pc54[18]);
FA1A GS54_19(ps55[18], pc55[19], g54[19], ps54[19], pc54[19]);
FA1A GS54_20(ps55[19], pc55[20], g54[20], ps54[20], pc54[20]);
FA1A GS54_21(ps55[20], pc55[21], g54[21], ps54[21], pc54[21]);
FA1A GS54_22(ps55[21], pc55[22], g54[22], ps54[22], pc54[22]);
FA1A GS54_23(ps55[22], pc55[23], g54[23], ps54[23], pc54[23]);
FA1A GS54_24(ps55[23], pc55[24], g54[24], ps54[24], pc54[24]);
FA1A GS54_25(ps55[24], pc55[25], g54[25], ps54[25], pc54[25]);
FA1A GS54_26(ps55[25], pc55[26], g54[26], ps54[26], pc54[26]);
FA1A GS54_27(ps55[26], pc55[27], g54[27], ps54[27], pc54[27]);
FA1A GS54_28(ps55[27], pc55[28], g54[28], ps54[28], pc54[28]);
FA1A GS54_29(ps55[28], pc55[29], g54[29], ps54[29], pc54[29]);
FA1A GS54_30(ps55[29], pc55[30], g54[30], ps54[30], pc54[30]);
FA1A GS54_31(ps55[30], pc55[31], g54[31], ps54[31], pc54[31]);
FA1A GS54_32(ps55[31], pc55[32], g54[32], ps54[32], pc54[32]);
FA1A GS54_33(ps55[32], pc55[33], g54[33], ps54[33], pc54[33]);
FA1A GS54_34(ps55[33], pc55[34], g54[34], ps54[34], pc54[34]);
FA1A GS54_35(ps55[34], pc55[35], g54[35], ps54[35], pc54[35]);
FA1A GS54_36(ps55[35], pc55[36], g54[36], ps54[36], pc54[36]);
FA1A GS54_37(ps55[36], pc55[37], g54[37], ps54[37], pc54[37]);
FA1A GS54_38(ps55[37], pc55[38], g54[38], ps54[38], pc54[38]);
FA1A GS54_39(ps55[38], pc55[39], g54[39], ps54[39], pc54[39]);
FA1A GS54_40(ps55[39], pc55[40], g54[40], ps54[40], pc54[40]);
FA1A GS54_41(ps55[40], pc55[41], g54[41], ps54[41], pc54[41]);
FA1A GS54_42(ps55[41], pc55[42], g54[42], ps54[42], pc54[42]);
FA1A GS54_43(ps55[42], pc55[43], g54[43], ps54[43], pc54[43]);
FA1A GS54_44(ps55[43], pc55[44], g54[44], ps54[44], pc54[44]);
FA1A GS54_45(ps55[44], pc55[45], g54[45], ps54[45], pc54[45]);
FA1A GS54_46(ps55[45], pc55[46], g54[46], ps54[46], pc54[46]);
FA1A GS54_47(ps55[46], pc55[47], g54[47], ps54[47], pc54[47]);
FA1A GS54_48(ps55[47], pc55[48], g54[48], ps54[48], pc54[48]);
FA1A GS54_49(ps55[48], pc55[49], g54[49], ps54[49], pc54[49]);
FA1A GS54_50(ps55[49], pc55[50], g54[50], ps54[50], pc54[50]);
FA1A GS54_51(ps55[50], pc55[51], g54[51], ps54[51], pc54[51]);
FA1A GS54_52(ps55[51], pc55[52], g54[52], ps54[52], pc54[52]);
FA1A GS54_53(ps55[52], pc55[53], g54[53], ps54[53], pc54[53]);
FA1A GS54_54(ps55[53], pc55[54], g54[54], ps54[54], pc54[54]);
FA1A GS54_55(ps55[54], pc55[55], g54[55], ps54[55], pc54[55]);
FA1A GS54_56(ps55[55], pc55[56], g54[56], ps54[56], pc54[56]);
FA1A GS54_57(ps55[56], pc55[57], g54[57], ps54[57], pc54[57]);
FA1A GS54_58(ps55[57], pc55[58], g54[58], ps54[58], pc54[58]);
FA1A GS54_59(ps55[58], pc55[59], g54[59], ps54[59], pc54[59]);
FA1A GS54_60(ps55[59], pc55[60], g54[60], ps54[60], pc54[60]);
FA1A GS54_61(ps55[60], pc55[61], g54[61], ps54[61], pc54[61]);
FA1A GS54_62(ps55[61], pc55[62], g54[62], ps54[62], pc54[62]);
FA1A GS54_63(ps55[62], pc55[63], g54[63], ps54[63], pc54[63]);
FA1A GS53_9(g54[8], pc54[9], g53[9], ps53[9], pc53[9]);
FA1A GS53_10(ps54[9], pc54[10], g53[10], ps53[10], pc53[10]);
FA1A GS53_11(ps54[10], pc54[11], g53[11], ps53[11], pc53[11]);
FA1A GS53_12(ps54[11], pc54[12], g53[12], ps53[12], pc53[12]);
FA1A GS53_13(ps54[12], pc54[13], g53[13], ps53[13], pc53[13]);
FA1A GS53_14(ps54[13], pc54[14], g53[14], ps53[14], pc53[14]);
FA1A GS53_15(ps54[14], pc54[15], g53[15], ps53[15], pc53[15]);
FA1A GS53_16(ps54[15], pc54[16], g53[16], ps53[16], pc53[16]);
FA1A GS53_17(ps54[16], pc54[17], g53[17], ps53[17], pc53[17]);
FA1A GS53_18(ps54[17], pc54[18], g53[18], ps53[18], pc53[18]);
FA1A GS53_19(ps54[18], pc54[19], g53[19], ps53[19], pc53[19]);
FA1A GS53_20(ps54[19], pc54[20], g53[20], ps53[20], pc53[20]);
FA1A GS53_21(ps54[20], pc54[21], g53[21], ps53[21], pc53[21]);
FA1A GS53_22(ps54[21], pc54[22], g53[22], ps53[22], pc53[22]);
FA1A GS53_23(ps54[22], pc54[23], g53[23], ps53[23], pc53[23]);
FA1A GS53_24(ps54[23], pc54[24], g53[24], ps53[24], pc53[24]);
FA1A GS53_25(ps54[24], pc54[25], g53[25], ps53[25], pc53[25]);
FA1A GS53_26(ps54[25], pc54[26], g53[26], ps53[26], pc53[26]);
FA1A GS53_27(ps54[26], pc54[27], g53[27], ps53[27], pc53[27]);
FA1A GS53_28(ps54[27], pc54[28], g53[28], ps53[28], pc53[28]);
FA1A GS53_29(ps54[28], pc54[29], g53[29], ps53[29], pc53[29]);
FA1A GS53_30(ps54[29], pc54[30], g53[30], ps53[30], pc53[30]);
FA1A GS53_31(ps54[30], pc54[31], g53[31], ps53[31], pc53[31]);
FA1A GS53_32(ps54[31], pc54[32], g53[32], ps53[32], pc53[32]);
FA1A GS53_33(ps54[32], pc54[33], g53[33], ps53[33], pc53[33]);
FA1A GS53_34(ps54[33], pc54[34], g53[34], ps53[34], pc53[34]);
FA1A GS53_35(ps54[34], pc54[35], g53[35], ps53[35], pc53[35]);
FA1A GS53_36(ps54[35], pc54[36], g53[36], ps53[36], pc53[36]);
FA1A GS53_37(ps54[36], pc54[37], g53[37], ps53[37], pc53[37]);
FA1A GS53_38(ps54[37], pc54[38], g53[38], ps53[38], pc53[38]);
FA1A GS53_39(ps54[38], pc54[39], g53[39], ps53[39], pc53[39]);
FA1A GS53_40(ps54[39], pc54[40], g53[40], ps53[40], pc53[40]);
FA1A GS53_41(ps54[40], pc54[41], g53[41], ps53[41], pc53[41]);
FA1A GS53_42(ps54[41], pc54[42], g53[42], ps53[42], pc53[42]);
FA1A GS53_43(ps54[42], pc54[43], g53[43], ps53[43], pc53[43]);
FA1A GS53_44(ps54[43], pc54[44], g53[44], ps53[44], pc53[44]);
FA1A GS53_45(ps54[44], pc54[45], g53[45], ps53[45], pc53[45]);
FA1A GS53_46(ps54[45], pc54[46], g53[46], ps53[46], pc53[46]);
FA1A GS53_47(ps54[46], pc54[47], g53[47], ps53[47], pc53[47]);
FA1A GS53_48(ps54[47], pc54[48], g53[48], ps53[48], pc53[48]);
FA1A GS53_49(ps54[48], pc54[49], g53[49], ps53[49], pc53[49]);
FA1A GS53_50(ps54[49], pc54[50], g53[50], ps53[50], pc53[50]);
FA1A GS53_51(ps54[50], pc54[51], g53[51], ps53[51], pc53[51]);
FA1A GS53_52(ps54[51], pc54[52], g53[52], ps53[52], pc53[52]);
FA1A GS53_53(ps54[52], pc54[53], g53[53], ps53[53], pc53[53]);
FA1A GS53_54(ps54[53], pc54[54], g53[54], ps53[54], pc53[54]);
FA1A GS53_55(ps54[54], pc54[55], g53[55], ps53[55], pc53[55]);
FA1A GS53_56(ps54[55], pc54[56], g53[56], ps53[56], pc53[56]);
FA1A GS53_57(ps54[56], pc54[57], g53[57], ps53[57], pc53[57]);
FA1A GS53_58(ps54[57], pc54[58], g53[58], ps53[58], pc53[58]);
FA1A GS53_59(ps54[58], pc54[59], g53[59], ps53[59], pc53[59]);
FA1A GS53_60(ps54[59], pc54[60], g53[60], ps53[60], pc53[60]);
FA1A GS53_61(ps54[60], pc54[61], g53[61], ps53[61], pc53[61]);
FA1A GS53_62(ps54[61], pc54[62], g53[62], ps53[62], pc53[62]);
FA1A GS53_63(ps54[62], pc54[63], g53[63], ps53[63], pc53[63]);
FA1A GS52_9(g53[8], pc53[9], g52[9], ps52[9], pc52[9]);
FA1A GS52_10(ps53[9], pc53[10], g52[10], ps52[10], pc52[10]);
FA1A GS52_11(ps53[10], pc53[11], g52[11], ps52[11], pc52[11]);
FA1A GS52_12(ps53[11], pc53[12], g52[12], ps52[12], pc52[12]);
FA1A GS52_13(ps53[12], pc53[13], g52[13], ps52[13], pc52[13]);
FA1A GS52_14(ps53[13], pc53[14], g52[14], ps52[14], pc52[14]);
FA1A GS52_15(ps53[14], pc53[15], g52[15], ps52[15], pc52[15]);
FA1A GS52_16(ps53[15], pc53[16], g52[16], ps52[16], pc52[16]);
FA1A GS52_17(ps53[16], pc53[17], g52[17], ps52[17], pc52[17]);
FA1A GS52_18(ps53[17], pc53[18], g52[18], ps52[18], pc52[18]);
FA1A GS52_19(ps53[18], pc53[19], g52[19], ps52[19], pc52[19]);
FA1A GS52_20(ps53[19], pc53[20], g52[20], ps52[20], pc52[20]);
FA1A GS52_21(ps53[20], pc53[21], g52[21], ps52[21], pc52[21]);
FA1A GS52_22(ps53[21], pc53[22], g52[22], ps52[22], pc52[22]);
FA1A GS52_23(ps53[22], pc53[23], g52[23], ps52[23], pc52[23]);
FA1A GS52_24(ps53[23], pc53[24], g52[24], ps52[24], pc52[24]);
FA1A GS52_25(ps53[24], pc53[25], g52[25], ps52[25], pc52[25]);
FA1A GS52_26(ps53[25], pc53[26], g52[26], ps52[26], pc52[26]);
FA1A GS52_27(ps53[26], pc53[27], g52[27], ps52[27], pc52[27]);
FA1A GS52_28(ps53[27], pc53[28], g52[28], ps52[28], pc52[28]);
FA1A GS52_29(ps53[28], pc53[29], g52[29], ps52[29], pc52[29]);
FA1A GS52_30(ps53[29], pc53[30], g52[30], ps52[30], pc52[30]);
FA1A GS52_31(ps53[30], pc53[31], g52[31], ps52[31], pc52[31]);
FA1A GS52_32(ps53[31], pc53[32], g52[32], ps52[32], pc52[32]);
FA1A GS52_33(ps53[32], pc53[33], g52[33], ps52[33], pc52[33]);
FA1A GS52_34(ps53[33], pc53[34], g52[34], ps52[34], pc52[34]);
FA1A GS52_35(ps53[34], pc53[35], g52[35], ps52[35], pc52[35]);
FA1A GS52_36(ps53[35], pc53[36], g52[36], ps52[36], pc52[36]);
FA1A GS52_37(ps53[36], pc53[37], g52[37], ps52[37], pc52[37]);
FA1A GS52_38(ps53[37], pc53[38], g52[38], ps52[38], pc52[38]);
FA1A GS52_39(ps53[38], pc53[39], g52[39], ps52[39], pc52[39]);
FA1A GS52_40(ps53[39], pc53[40], g52[40], ps52[40], pc52[40]);
FA1A GS52_41(ps53[40], pc53[41], g52[41], ps52[41], pc52[41]);
FA1A GS52_42(ps53[41], pc53[42], g52[42], ps52[42], pc52[42]);
FA1A GS52_43(ps53[42], pc53[43], g52[43], ps52[43], pc52[43]);
FA1A GS52_44(ps53[43], pc53[44], g52[44], ps52[44], pc52[44]);
FA1A GS52_45(ps53[44], pc53[45], g52[45], ps52[45], pc52[45]);
FA1A GS52_46(ps53[45], pc53[46], g52[46], ps52[46], pc52[46]);
FA1A GS52_47(ps53[46], pc53[47], g52[47], ps52[47], pc52[47]);
FA1A GS52_48(ps53[47], pc53[48], g52[48], ps52[48], pc52[48]);
FA1A GS52_49(ps53[48], pc53[49], g52[49], ps52[49], pc52[49]);
FA1A GS52_50(ps53[49], pc53[50], g52[50], ps52[50], pc52[50]);
FA1A GS52_51(ps53[50], pc53[51], g52[51], ps52[51], pc52[51]);
FA1A GS52_52(ps53[51], pc53[52], g52[52], ps52[52], pc52[52]);
FA1A GS52_53(ps53[52], pc53[53], g52[53], ps52[53], pc52[53]);
FA1A GS52_54(ps53[53], pc53[54], g52[54], ps52[54], pc52[54]);
FA1A GS52_55(ps53[54], pc53[55], g52[55], ps52[55], pc52[55]);
FA1A GS52_56(ps53[55], pc53[56], g52[56], ps52[56], pc52[56]);
FA1A GS52_57(ps53[56], pc53[57], g52[57], ps52[57], pc52[57]);
FA1A GS52_58(ps53[57], pc53[58], g52[58], ps52[58], pc52[58]);
FA1A GS52_59(ps53[58], pc53[59], g52[59], ps52[59], pc52[59]);
FA1A GS52_60(ps53[59], pc53[60], g52[60], ps52[60], pc52[60]);
FA1A GS52_61(ps53[60], pc53[61], g52[61], ps52[61], pc52[61]);
FA1A GS52_62(ps53[61], pc53[62], g52[62], ps52[62], pc52[62]);
FA1A GS52_63(ps53[62], pc53[63], g52[63], ps52[63], pc52[63]);
FA1A GS51_9(g52[8], pc52[9], g51[9], ps51[9], pc51[9]);
FA1A GS51_10(ps52[9], pc52[10], g51[10], ps51[10], pc51[10]);
FA1A GS51_11(ps52[10], pc52[11], g51[11], ps51[11], pc51[11]);
FA1A GS51_12(ps52[11], pc52[12], g51[12], ps51[12], pc51[12]);
FA1A GS51_13(ps52[12], pc52[13], g51[13], ps51[13], pc51[13]);
FA1A GS51_14(ps52[13], pc52[14], g51[14], ps51[14], pc51[14]);
FA1A GS51_15(ps52[14], pc52[15], g51[15], ps51[15], pc51[15]);
FA1A GS51_16(ps52[15], pc52[16], g51[16], ps51[16], pc51[16]);
FA1A GS51_17(ps52[16], pc52[17], g51[17], ps51[17], pc51[17]);
FA1A GS51_18(ps52[17], pc52[18], g51[18], ps51[18], pc51[18]);
FA1A GS51_19(ps52[18], pc52[19], g51[19], ps51[19], pc51[19]);
FA1A GS51_20(ps52[19], pc52[20], g51[20], ps51[20], pc51[20]);
FA1A GS51_21(ps52[20], pc52[21], g51[21], ps51[21], pc51[21]);
FA1A GS51_22(ps52[21], pc52[22], g51[22], ps51[22], pc51[22]);
FA1A GS51_23(ps52[22], pc52[23], g51[23], ps51[23], pc51[23]);
FA1A GS51_24(ps52[23], pc52[24], g51[24], ps51[24], pc51[24]);
FA1A GS51_25(ps52[24], pc52[25], g51[25], ps51[25], pc51[25]);
FA1A GS51_26(ps52[25], pc52[26], g51[26], ps51[26], pc51[26]);
FA1A GS51_27(ps52[26], pc52[27], g51[27], ps51[27], pc51[27]);
FA1A GS51_28(ps52[27], pc52[28], g51[28], ps51[28], pc51[28]);
FA1A GS51_29(ps52[28], pc52[29], g51[29], ps51[29], pc51[29]);
FA1A GS51_30(ps52[29], pc52[30], g51[30], ps51[30], pc51[30]);
FA1A GS51_31(ps52[30], pc52[31], g51[31], ps51[31], pc51[31]);
FA1A GS51_32(ps52[31], pc52[32], g51[32], ps51[32], pc51[32]);
FA1A GS51_33(ps52[32], pc52[33], g51[33], ps51[33], pc51[33]);
FA1A GS51_34(ps52[33], pc52[34], g51[34], ps51[34], pc51[34]);
FA1A GS51_35(ps52[34], pc52[35], g51[35], ps51[35], pc51[35]);
FA1A GS51_36(ps52[35], pc52[36], g51[36], ps51[36], pc51[36]);
FA1A GS51_37(ps52[36], pc52[37], g51[37], ps51[37], pc51[37]);
FA1A GS51_38(ps52[37], pc52[38], g51[38], ps51[38], pc51[38]);
FA1A GS51_39(ps52[38], pc52[39], g51[39], ps51[39], pc51[39]);
FA1A GS51_40(ps52[39], pc52[40], g51[40], ps51[40], pc51[40]);
FA1A GS51_41(ps52[40], pc52[41], g51[41], ps51[41], pc51[41]);
FA1A GS51_42(ps52[41], pc52[42], g51[42], ps51[42], pc51[42]);
FA1A GS51_43(ps52[42], pc52[43], g51[43], ps51[43], pc51[43]);
FA1A GS51_44(ps52[43], pc52[44], g51[44], ps51[44], pc51[44]);
FA1A GS51_45(ps52[44], pc52[45], g51[45], ps51[45], pc51[45]);
FA1A GS51_46(ps52[45], pc52[46], g51[46], ps51[46], pc51[46]);
FA1A GS51_47(ps52[46], pc52[47], g51[47], ps51[47], pc51[47]);
FA1A GS51_48(ps52[47], pc52[48], g51[48], ps51[48], pc51[48]);
FA1A GS51_49(ps52[48], pc52[49], g51[49], ps51[49], pc51[49]);
FA1A GS51_50(ps52[49], pc52[50], g51[50], ps51[50], pc51[50]);
FA1A GS51_51(ps52[50], pc52[51], g51[51], ps51[51], pc51[51]);
FA1A GS51_52(ps52[51], pc52[52], g51[52], ps51[52], pc51[52]);
FA1A GS51_53(ps52[52], pc52[53], g51[53], ps51[53], pc51[53]);
FA1A GS51_54(ps52[53], pc52[54], g51[54], ps51[54], pc51[54]);
FA1A GS51_55(ps52[54], pc52[55], g51[55], ps51[55], pc51[55]);
FA1A GS51_56(ps52[55], pc52[56], g51[56], ps51[56], pc51[56]);
FA1A GS51_57(ps52[56], pc52[57], g51[57], ps51[57], pc51[57]);
FA1A GS51_58(ps52[57], pc52[58], g51[58], ps51[58], pc51[58]);
FA1A GS51_59(ps52[58], pc52[59], g51[59], ps51[59], pc51[59]);
FA1A GS51_60(ps52[59], pc52[60], g51[60], ps51[60], pc51[60]);
FA1A GS51_61(ps52[60], pc52[61], g51[61], ps51[61], pc51[61]);
FA1A GS51_62(ps52[61], pc52[62], g51[62], ps51[62], pc51[62]);
FA1A GS51_63(ps52[62], pc52[63], g51[63], ps51[63], pc51[63]);
FA1A GS50_9(g51[8], pc51[9], g50[9], ps50[9], pc50[9]);
FA1A GS50_10(ps51[9], pc51[10], g50[10], ps50[10], pc50[10]);
FA1A GS50_11(ps51[10], pc51[11], g50[11], ps50[11], pc50[11]);
FA1A GS50_12(ps51[11], pc51[12], g50[12], ps50[12], pc50[12]);
FA1A GS50_13(ps51[12], pc51[13], g50[13], ps50[13], pc50[13]);
FA1A GS50_14(ps51[13], pc51[14], g50[14], ps50[14], pc50[14]);
FA1A GS50_15(ps51[14], pc51[15], g50[15], ps50[15], pc50[15]);
FA1A GS50_16(ps51[15], pc51[16], g50[16], ps50[16], pc50[16]);
FA1A GS50_17(ps51[16], pc51[17], g50[17], ps50[17], pc50[17]);
FA1A GS50_18(ps51[17], pc51[18], g50[18], ps50[18], pc50[18]);
FA1A GS50_19(ps51[18], pc51[19], g50[19], ps50[19], pc50[19]);
FA1A GS50_20(ps51[19], pc51[20], g50[20], ps50[20], pc50[20]);
FA1A GS50_21(ps51[20], pc51[21], g50[21], ps50[21], pc50[21]);
FA1A GS50_22(ps51[21], pc51[22], g50[22], ps50[22], pc50[22]);
FA1A GS50_23(ps51[22], pc51[23], g50[23], ps50[23], pc50[23]);
FA1A GS50_24(ps51[23], pc51[24], g50[24], ps50[24], pc50[24]);
FA1A GS50_25(ps51[24], pc51[25], g50[25], ps50[25], pc50[25]);
FA1A GS50_26(ps51[25], pc51[26], g50[26], ps50[26], pc50[26]);
FA1A GS50_27(ps51[26], pc51[27], g50[27], ps50[27], pc50[27]);
FA1A GS50_28(ps51[27], pc51[28], g50[28], ps50[28], pc50[28]);
FA1A GS50_29(ps51[28], pc51[29], g50[29], ps50[29], pc50[29]);
FA1A GS50_30(ps51[29], pc51[30], g50[30], ps50[30], pc50[30]);
FA1A GS50_31(ps51[30], pc51[31], g50[31], ps50[31], pc50[31]);
FA1A GS50_32(ps51[31], pc51[32], g50[32], ps50[32], pc50[32]);
FA1A GS50_33(ps51[32], pc51[33], g50[33], ps50[33], pc50[33]);
FA1A GS50_34(ps51[33], pc51[34], g50[34], ps50[34], pc50[34]);
FA1A GS50_35(ps51[34], pc51[35], g50[35], ps50[35], pc50[35]);
FA1A GS50_36(ps51[35], pc51[36], g50[36], ps50[36], pc50[36]);
FA1A GS50_37(ps51[36], pc51[37], g50[37], ps50[37], pc50[37]);
FA1A GS50_38(ps51[37], pc51[38], g50[38], ps50[38], pc50[38]);
FA1A GS50_39(ps51[38], pc51[39], g50[39], ps50[39], pc50[39]);
FA1A GS50_40(ps51[39], pc51[40], g50[40], ps50[40], pc50[40]);
FA1A GS50_41(ps51[40], pc51[41], g50[41], ps50[41], pc50[41]);
FA1A GS50_42(ps51[41], pc51[42], g50[42], ps50[42], pc50[42]);
FA1A GS50_43(ps51[42], pc51[43], g50[43], ps50[43], pc50[43]);
FA1A GS50_44(ps51[43], pc51[44], g50[44], ps50[44], pc50[44]);
FA1A GS50_45(ps51[44], pc51[45], g50[45], ps50[45], pc50[45]);
FA1A GS50_46(ps51[45], pc51[46], g50[46], ps50[46], pc50[46]);
FA1A GS50_47(ps51[46], pc51[47], g50[47], ps50[47], pc50[47]);
FA1A GS50_48(ps51[47], pc51[48], g50[48], ps50[48], pc50[48]);
FA1A GS50_49(ps51[48], pc51[49], g50[49], ps50[49], pc50[49]);
FA1A GS50_50(ps51[49], pc51[50], g50[50], ps50[50], pc50[50]);
FA1A GS50_51(ps51[50], pc51[51], g50[51], ps50[51], pc50[51]);
FA1A GS50_52(ps51[51], pc51[52], g50[52], ps50[52], pc50[52]);
FA1A GS50_53(ps51[52], pc51[53], g50[53], ps50[53], pc50[53]);
FA1A GS50_54(ps51[53], pc51[54], g50[54], ps50[54], pc50[54]);
FA1A GS50_55(ps51[54], pc51[55], g50[55], ps50[55], pc50[55]);
FA1A GS50_56(ps51[55], pc51[56], g50[56], ps50[56], pc50[56]);
FA1A GS50_57(ps51[56], pc51[57], g50[57], ps50[57], pc50[57]);
FA1A GS50_58(ps51[57], pc51[58], g50[58], ps50[58], pc50[58]);
FA1A GS50_59(ps51[58], pc51[59], g50[59], ps50[59], pc50[59]);
FA1A GS50_60(ps51[59], pc51[60], g50[60], ps50[60], pc50[60]);
FA1A GS50_61(ps51[60], pc51[61], g50[61], ps50[61], pc50[61]);
FA1A GS50_62(ps51[61], pc51[62], g50[62], ps50[62], pc50[62]);
FA1A GS50_63(ps51[62], pc51[63], g50[63], ps50[63], pc50[63]);
FA1A GS49_9(g50[8], pc50[9], g49[9], ps49[9], pc49[9]);
FA1A GS49_10(ps50[9], pc50[10], g49[10], ps49[10], pc49[10]);
FA1A GS49_11(ps50[10], pc50[11], g49[11], ps49[11], pc49[11]);
FA1A GS49_12(ps50[11], pc50[12], g49[12], ps49[12], pc49[12]);
FA1A GS49_13(ps50[12], pc50[13], g49[13], ps49[13], pc49[13]);
FA1A GS49_14(ps50[13], pc50[14], g49[14], ps49[14], pc49[14]);
FA1A GS49_15(ps50[14], pc50[15], g49[15], ps49[15], pc49[15]);
FA1A GS49_16(ps50[15], pc50[16], g49[16], ps49[16], pc49[16]);
FA1A GS49_17(ps50[16], pc50[17], g49[17], ps49[17], pc49[17]);
FA1A GS49_18(ps50[17], pc50[18], g49[18], ps49[18], pc49[18]);
FA1A GS49_19(ps50[18], pc50[19], g49[19], ps49[19], pc49[19]);
FA1A GS49_20(ps50[19], pc50[20], g49[20], ps49[20], pc49[20]);
FA1A GS49_21(ps50[20], pc50[21], g49[21], ps49[21], pc49[21]);
FA1A GS49_22(ps50[21], pc50[22], g49[22], ps49[22], pc49[22]);
FA1A GS49_23(ps50[22], pc50[23], g49[23], ps49[23], pc49[23]);
FA1A GS49_24(ps50[23], pc50[24], g49[24], ps49[24], pc49[24]);
FA1A GS49_25(ps50[24], pc50[25], g49[25], ps49[25], pc49[25]);
FA1A GS49_26(ps50[25], pc50[26], g49[26], ps49[26], pc49[26]);
FA1A GS49_27(ps50[26], pc50[27], g49[27], ps49[27], pc49[27]);
FA1A GS49_28(ps50[27], pc50[28], g49[28], ps49[28], pc49[28]);
FA1A GS49_29(ps50[28], pc50[29], g49[29], ps49[29], pc49[29]);
FA1A GS49_30(ps50[29], pc50[30], g49[30], ps49[30], pc49[30]);
FA1A GS49_31(ps50[30], pc50[31], g49[31], ps49[31], pc49[31]);
FA1A GS49_32(ps50[31], pc50[32], g49[32], ps49[32], pc49[32]);
FA1A GS49_33(ps50[32], pc50[33], g49[33], ps49[33], pc49[33]);
FA1A GS49_34(ps50[33], pc50[34], g49[34], ps49[34], pc49[34]);
FA1A GS49_35(ps50[34], pc50[35], g49[35], ps49[35], pc49[35]);
FA1A GS49_36(ps50[35], pc50[36], g49[36], ps49[36], pc49[36]);
FA1A GS49_37(ps50[36], pc50[37], g49[37], ps49[37], pc49[37]);
FA1A GS49_38(ps50[37], pc50[38], g49[38], ps49[38], pc49[38]);
FA1A GS49_39(ps50[38], pc50[39], g49[39], ps49[39], pc49[39]);
FA1A GS49_40(ps50[39], pc50[40], g49[40], ps49[40], pc49[40]);
FA1A GS49_41(ps50[40], pc50[41], g49[41], ps49[41], pc49[41]);
FA1A GS49_42(ps50[41], pc50[42], g49[42], ps49[42], pc49[42]);
FA1A GS49_43(ps50[42], pc50[43], g49[43], ps49[43], pc49[43]);
FA1A GS49_44(ps50[43], pc50[44], g49[44], ps49[44], pc49[44]);
FA1A GS49_45(ps50[44], pc50[45], g49[45], ps49[45], pc49[45]);
FA1A GS49_46(ps50[45], pc50[46], g49[46], ps49[46], pc49[46]);
FA1A GS49_47(ps50[46], pc50[47], g49[47], ps49[47], pc49[47]);
FA1A GS49_48(ps50[47], pc50[48], g49[48], ps49[48], pc49[48]);
FA1A GS49_49(ps50[48], pc50[49], g49[49], ps49[49], pc49[49]);
FA1A GS49_50(ps50[49], pc50[50], g49[50], ps49[50], pc49[50]);
FA1A GS49_51(ps50[50], pc50[51], g49[51], ps49[51], pc49[51]);
FA1A GS49_52(ps50[51], pc50[52], g49[52], ps49[52], pc49[52]);
FA1A GS49_53(ps50[52], pc50[53], g49[53], ps49[53], pc49[53]);
FA1A GS49_54(ps50[53], pc50[54], g49[54], ps49[54], pc49[54]);
FA1A GS49_55(ps50[54], pc50[55], g49[55], ps49[55], pc49[55]);
FA1A GS49_56(ps50[55], pc50[56], g49[56], ps49[56], pc49[56]);
FA1A GS49_57(ps50[56], pc50[57], g49[57], ps49[57], pc49[57]);
FA1A GS49_58(ps50[57], pc50[58], g49[58], ps49[58], pc49[58]);
FA1A GS49_59(ps50[58], pc50[59], g49[59], ps49[59], pc49[59]);
FA1A GS49_60(ps50[59], pc50[60], g49[60], ps49[60], pc49[60]);
FA1A GS49_61(ps50[60], pc50[61], g49[61], ps49[61], pc49[61]);
FA1A GS49_62(ps50[61], pc50[62], g49[62], ps49[62], pc49[62]);
FA1A GS49_63(ps50[62], pc50[63], g49[63], ps49[63], pc49[63]);
FA1A GS48_9(g49[8], pc49[9], g48[9], ps48[9], pc48[9]);
FA1A GS48_10(ps49[9], pc49[10], g48[10], ps48[10], pc48[10]);
FA1A GS48_11(ps49[10], pc49[11], g48[11], ps48[11], pc48[11]);
FA1A GS48_12(ps49[11], pc49[12], g48[12], ps48[12], pc48[12]);
FA1A GS48_13(ps49[12], pc49[13], g48[13], ps48[13], pc48[13]);
FA1A GS48_14(ps49[13], pc49[14], g48[14], ps48[14], pc48[14]);
FA1A GS48_15(ps49[14], pc49[15], g48[15], ps48[15], pc48[15]);
FA1A GS48_16(ps49[15], pc49[16], g48[16], ps48[16], pc48[16]);
FA1A GS48_17(ps49[16], pc49[17], g48[17], ps48[17], pc48[17]);
FA1A GS48_18(ps49[17], pc49[18], g48[18], ps48[18], pc48[18]);
FA1A GS48_19(ps49[18], pc49[19], g48[19], ps48[19], pc48[19]);
FA1A GS48_20(ps49[19], pc49[20], g48[20], ps48[20], pc48[20]);
FA1A GS48_21(ps49[20], pc49[21], g48[21], ps48[21], pc48[21]);
FA1A GS48_22(ps49[21], pc49[22], g48[22], ps48[22], pc48[22]);
FA1A GS48_23(ps49[22], pc49[23], g48[23], ps48[23], pc48[23]);
FA1A GS48_24(ps49[23], pc49[24], g48[24], ps48[24], pc48[24]);
FA1A GS48_25(ps49[24], pc49[25], g48[25], ps48[25], pc48[25]);
FA1A GS48_26(ps49[25], pc49[26], g48[26], ps48[26], pc48[26]);
FA1A GS48_27(ps49[26], pc49[27], g48[27], ps48[27], pc48[27]);
FA1A GS48_28(ps49[27], pc49[28], g48[28], ps48[28], pc48[28]);
FA1A GS48_29(ps49[28], pc49[29], g48[29], ps48[29], pc48[29]);
FA1A GS48_30(ps49[29], pc49[30], g48[30], ps48[30], pc48[30]);
FA1A GS48_31(ps49[30], pc49[31], g48[31], ps48[31], pc48[31]);
FA1A GS48_32(ps49[31], pc49[32], g48[32], ps48[32], pc48[32]);
FA1A GS48_33(ps49[32], pc49[33], g48[33], ps48[33], pc48[33]);
FA1A GS48_34(ps49[33], pc49[34], g48[34], ps48[34], pc48[34]);
FA1A GS48_35(ps49[34], pc49[35], g48[35], ps48[35], pc48[35]);
FA1A GS48_36(ps49[35], pc49[36], g48[36], ps48[36], pc48[36]);
FA1A GS48_37(ps49[36], pc49[37], g48[37], ps48[37], pc48[37]);
FA1A GS48_38(ps49[37], pc49[38], g48[38], ps48[38], pc48[38]);
FA1A GS48_39(ps49[38], pc49[39], g48[39], ps48[39], pc48[39]);
FA1A GS48_40(ps49[39], pc49[40], g48[40], ps48[40], pc48[40]);
FA1A GS48_41(ps49[40], pc49[41], g48[41], ps48[41], pc48[41]);
FA1A GS48_42(ps49[41], pc49[42], g48[42], ps48[42], pc48[42]);
FA1A GS48_43(ps49[42], pc49[43], g48[43], ps48[43], pc48[43]);
FA1A GS48_44(ps49[43], pc49[44], g48[44], ps48[44], pc48[44]);
FA1A GS48_45(ps49[44], pc49[45], g48[45], ps48[45], pc48[45]);
FA1A GS48_46(ps49[45], pc49[46], g48[46], ps48[46], pc48[46]);
FA1A GS48_47(ps49[46], pc49[47], g48[47], ps48[47], pc48[47]);
FA1A GS48_48(ps49[47], pc49[48], g48[48], ps48[48], pc48[48]);
FA1A GS48_49(ps49[48], pc49[49], g48[49], ps48[49], pc48[49]);
FA1A GS48_50(ps49[49], pc49[50], g48[50], ps48[50], pc48[50]);
FA1A GS48_51(ps49[50], pc49[51], g48[51], ps48[51], pc48[51]);
FA1A GS48_52(ps49[51], pc49[52], g48[52], ps48[52], pc48[52]);
FA1A GS48_53(ps49[52], pc49[53], g48[53], ps48[53], pc48[53]);
FA1A GS48_54(ps49[53], pc49[54], g48[54], ps48[54], pc48[54]);
FA1A GS48_55(ps49[54], pc49[55], g48[55], ps48[55], pc48[55]);
FA1A GS48_56(ps49[55], pc49[56], g48[56], ps48[56], pc48[56]);
FA1A GS48_57(ps49[56], pc49[57], g48[57], ps48[57], pc48[57]);
FA1A GS48_58(ps49[57], pc49[58], g48[58], ps48[58], pc48[58]);
FA1A GS48_59(ps49[58], pc49[59], g48[59], ps48[59], pc48[59]);
FA1A GS48_60(ps49[59], pc49[60], g48[60], ps48[60], pc48[60]);
FA1A GS48_61(ps49[60], pc49[61], g48[61], ps48[61], pc48[61]);
FA1A GS48_62(ps49[61], pc49[62], g48[62], ps48[62], pc48[62]);
FA1A GS48_63(ps49[62], pc49[63], g48[63], ps48[63], pc48[63]);
FA1A GS47_9(g48[8], pc48[9], g47[9], ps47[9], pc47[9]);
FA1A GS47_10(ps48[9], pc48[10], g47[10], ps47[10], pc47[10]);
FA1A GS47_11(ps48[10], pc48[11], g47[11], ps47[11], pc47[11]);
FA1A GS47_12(ps48[11], pc48[12], g47[12], ps47[12], pc47[12]);
FA1A GS47_13(ps48[12], pc48[13], g47[13], ps47[13], pc47[13]);
FA1A GS47_14(ps48[13], pc48[14], g47[14], ps47[14], pc47[14]);
FA1A GS47_15(ps48[14], pc48[15], g47[15], ps47[15], pc47[15]);
FA1A GS47_16(ps48[15], pc48[16], g47[16], ps47[16], pc47[16]);
FA1A GS47_17(ps48[16], pc48[17], g47[17], ps47[17], pc47[17]);
FA1A GS47_18(ps48[17], pc48[18], g47[18], ps47[18], pc47[18]);
FA1A GS47_19(ps48[18], pc48[19], g47[19], ps47[19], pc47[19]);
FA1A GS47_20(ps48[19], pc48[20], g47[20], ps47[20], pc47[20]);
FA1A GS47_21(ps48[20], pc48[21], g47[21], ps47[21], pc47[21]);
FA1A GS47_22(ps48[21], pc48[22], g47[22], ps47[22], pc47[22]);
FA1A GS47_23(ps48[22], pc48[23], g47[23], ps47[23], pc47[23]);
FA1A GS47_24(ps48[23], pc48[24], g47[24], ps47[24], pc47[24]);
FA1A GS47_25(ps48[24], pc48[25], g47[25], ps47[25], pc47[25]);
FA1A GS47_26(ps48[25], pc48[26], g47[26], ps47[26], pc47[26]);
FA1A GS47_27(ps48[26], pc48[27], g47[27], ps47[27], pc47[27]);
FA1A GS47_28(ps48[27], pc48[28], g47[28], ps47[28], pc47[28]);
FA1A GS47_29(ps48[28], pc48[29], g47[29], ps47[29], pc47[29]);
FA1A GS47_30(ps48[29], pc48[30], g47[30], ps47[30], pc47[30]);
FA1A GS47_31(ps48[30], pc48[31], g47[31], ps47[31], pc47[31]);
FA1A GS47_32(ps48[31], pc48[32], g47[32], ps47[32], pc47[32]);
FA1A GS47_33(ps48[32], pc48[33], g47[33], ps47[33], pc47[33]);
FA1A GS47_34(ps48[33], pc48[34], g47[34], ps47[34], pc47[34]);
FA1A GS47_35(ps48[34], pc48[35], g47[35], ps47[35], pc47[35]);
FA1A GS47_36(ps48[35], pc48[36], g47[36], ps47[36], pc47[36]);
FA1A GS47_37(ps48[36], pc48[37], g47[37], ps47[37], pc47[37]);
FA1A GS47_38(ps48[37], pc48[38], g47[38], ps47[38], pc47[38]);
FA1A GS47_39(ps48[38], pc48[39], g47[39], ps47[39], pc47[39]);
FA1A GS47_40(ps48[39], pc48[40], g47[40], ps47[40], pc47[40]);
FA1A GS47_41(ps48[40], pc48[41], g47[41], ps47[41], pc47[41]);
FA1A GS47_42(ps48[41], pc48[42], g47[42], ps47[42], pc47[42]);
FA1A GS47_43(ps48[42], pc48[43], g47[43], ps47[43], pc47[43]);
FA1A GS47_44(ps48[43], pc48[44], g47[44], ps47[44], pc47[44]);
FA1A GS47_45(ps48[44], pc48[45], g47[45], ps47[45], pc47[45]);
FA1A GS47_46(ps48[45], pc48[46], g47[46], ps47[46], pc47[46]);
FA1A GS47_47(ps48[46], pc48[47], g47[47], ps47[47], pc47[47]);
FA1A GS47_48(ps48[47], pc48[48], g47[48], ps47[48], pc47[48]);
FA1A GS47_49(ps48[48], pc48[49], g47[49], ps47[49], pc47[49]);
FA1A GS47_50(ps48[49], pc48[50], g47[50], ps47[50], pc47[50]);
FA1A GS47_51(ps48[50], pc48[51], g47[51], ps47[51], pc47[51]);
FA1A GS47_52(ps48[51], pc48[52], g47[52], ps47[52], pc47[52]);
FA1A GS47_53(ps48[52], pc48[53], g47[53], ps47[53], pc47[53]);
FA1A GS47_54(ps48[53], pc48[54], g47[54], ps47[54], pc47[54]);
FA1A GS47_55(ps48[54], pc48[55], g47[55], ps47[55], pc47[55]);
FA1A GS47_56(ps48[55], pc48[56], g47[56], ps47[56], pc47[56]);
FA1A GS47_57(ps48[56], pc48[57], g47[57], ps47[57], pc47[57]);
FA1A GS47_58(ps48[57], pc48[58], g47[58], ps47[58], pc47[58]);
FA1A GS47_59(ps48[58], pc48[59], g47[59], ps47[59], pc47[59]);
FA1A GS47_60(ps48[59], pc48[60], g47[60], ps47[60], pc47[60]);
FA1A GS47_61(ps48[60], pc48[61], g47[61], ps47[61], pc47[61]);
FA1A GS47_62(ps48[61], pc48[62], g47[62], ps47[62], pc47[62]);
FA1A GS47_63(ps48[62], pc48[63], g47[63], ps47[63], pc47[63]);
FA1A GS46_9(g47[8], pc47[9], g46[9], ps46[9], pc46[9]);
FA1A GS46_10(ps47[9], pc47[10], g46[10], ps46[10], pc46[10]);
FA1A GS46_11(ps47[10], pc47[11], g46[11], ps46[11], pc46[11]);
FA1A GS46_12(ps47[11], pc47[12], g46[12], ps46[12], pc46[12]);
FA1A GS46_13(ps47[12], pc47[13], g46[13], ps46[13], pc46[13]);
FA1A GS46_14(ps47[13], pc47[14], g46[14], ps46[14], pc46[14]);
FA1A GS46_15(ps47[14], pc47[15], g46[15], ps46[15], pc46[15]);
FA1A GS46_16(ps47[15], pc47[16], g46[16], ps46[16], pc46[16]);
FA1A GS46_17(ps47[16], pc47[17], g46[17], ps46[17], pc46[17]);
FA1A GS46_18(ps47[17], pc47[18], g46[18], ps46[18], pc46[18]);
FA1A GS46_19(ps47[18], pc47[19], g46[19], ps46[19], pc46[19]);
FA1A GS46_20(ps47[19], pc47[20], g46[20], ps46[20], pc46[20]);
FA1A GS46_21(ps47[20], pc47[21], g46[21], ps46[21], pc46[21]);
FA1A GS46_22(ps47[21], pc47[22], g46[22], ps46[22], pc46[22]);
FA1A GS46_23(ps47[22], pc47[23], g46[23], ps46[23], pc46[23]);
FA1A GS46_24(ps47[23], pc47[24], g46[24], ps46[24], pc46[24]);
FA1A GS46_25(ps47[24], pc47[25], g46[25], ps46[25], pc46[25]);
FA1A GS46_26(ps47[25], pc47[26], g46[26], ps46[26], pc46[26]);
FA1A GS46_27(ps47[26], pc47[27], g46[27], ps46[27], pc46[27]);
FA1A GS46_28(ps47[27], pc47[28], g46[28], ps46[28], pc46[28]);
FA1A GS46_29(ps47[28], pc47[29], g46[29], ps46[29], pc46[29]);
FA1A GS46_30(ps47[29], pc47[30], g46[30], ps46[30], pc46[30]);
FA1A GS46_31(ps47[30], pc47[31], g46[31], ps46[31], pc46[31]);
FA1A GS46_32(ps47[31], pc47[32], g46[32], ps46[32], pc46[32]);
FA1A GS46_33(ps47[32], pc47[33], g46[33], ps46[33], pc46[33]);
FA1A GS46_34(ps47[33], pc47[34], g46[34], ps46[34], pc46[34]);
FA1A GS46_35(ps47[34], pc47[35], g46[35], ps46[35], pc46[35]);
FA1A GS46_36(ps47[35], pc47[36], g46[36], ps46[36], pc46[36]);
FA1A GS46_37(ps47[36], pc47[37], g46[37], ps46[37], pc46[37]);
FA1A GS46_38(ps47[37], pc47[38], g46[38], ps46[38], pc46[38]);
FA1A GS46_39(ps47[38], pc47[39], g46[39], ps46[39], pc46[39]);
FA1A GS46_40(ps47[39], pc47[40], g46[40], ps46[40], pc46[40]);
FA1A GS46_41(ps47[40], pc47[41], g46[41], ps46[41], pc46[41]);
FA1A GS46_42(ps47[41], pc47[42], g46[42], ps46[42], pc46[42]);
FA1A GS46_43(ps47[42], pc47[43], g46[43], ps46[43], pc46[43]);
FA1A GS46_44(ps47[43], pc47[44], g46[44], ps46[44], pc46[44]);
FA1A GS46_45(ps47[44], pc47[45], g46[45], ps46[45], pc46[45]);
FA1A GS46_46(ps47[45], pc47[46], g46[46], ps46[46], pc46[46]);
FA1A GS46_47(ps47[46], pc47[47], g46[47], ps46[47], pc46[47]);
FA1A GS46_48(ps47[47], pc47[48], g46[48], ps46[48], pc46[48]);
FA1A GS46_49(ps47[48], pc47[49], g46[49], ps46[49], pc46[49]);
FA1A GS46_50(ps47[49], pc47[50], g46[50], ps46[50], pc46[50]);
FA1A GS46_51(ps47[50], pc47[51], g46[51], ps46[51], pc46[51]);
FA1A GS46_52(ps47[51], pc47[52], g46[52], ps46[52], pc46[52]);
FA1A GS46_53(ps47[52], pc47[53], g46[53], ps46[53], pc46[53]);
FA1A GS46_54(ps47[53], pc47[54], g46[54], ps46[54], pc46[54]);
FA1A GS46_55(ps47[54], pc47[55], g46[55], ps46[55], pc46[55]);
FA1A GS46_56(ps47[55], pc47[56], g46[56], ps46[56], pc46[56]);
FA1A GS46_57(ps47[56], pc47[57], g46[57], ps46[57], pc46[57]);
FA1A GS46_58(ps47[57], pc47[58], g46[58], ps46[58], pc46[58]);
FA1A GS46_59(ps47[58], pc47[59], g46[59], ps46[59], pc46[59]);
FA1A GS46_60(ps47[59], pc47[60], g46[60], ps46[60], pc46[60]);
FA1A GS46_61(ps47[60], pc47[61], g46[61], ps46[61], pc46[61]);
FA1A GS46_62(ps47[61], pc47[62], g46[62], ps46[62], pc46[62]);
FA1A GS46_63(ps47[62], pc47[63], g46[63], ps46[63], pc46[63]);
FA1A GS45_9(g46[8], pc46[9], g45[9], ps45[9], pc45[9]);
FA1A GS45_10(ps46[9], pc46[10], g45[10], ps45[10], pc45[10]);
FA1A GS45_11(ps46[10], pc46[11], g45[11], ps45[11], pc45[11]);
FA1A GS45_12(ps46[11], pc46[12], g45[12], ps45[12], pc45[12]);
FA1A GS45_13(ps46[12], pc46[13], g45[13], ps45[13], pc45[13]);
FA1A GS45_14(ps46[13], pc46[14], g45[14], ps45[14], pc45[14]);
FA1A GS45_15(ps46[14], pc46[15], g45[15], ps45[15], pc45[15]);
FA1A GS45_16(ps46[15], pc46[16], g45[16], ps45[16], pc45[16]);
FA1A GS45_17(ps46[16], pc46[17], g45[17], ps45[17], pc45[17]);
FA1A GS45_18(ps46[17], pc46[18], g45[18], ps45[18], pc45[18]);
FA1A GS45_19(ps46[18], pc46[19], g45[19], ps45[19], pc45[19]);
FA1A GS45_20(ps46[19], pc46[20], g45[20], ps45[20], pc45[20]);
FA1A GS45_21(ps46[20], pc46[21], g45[21], ps45[21], pc45[21]);
FA1A GS45_22(ps46[21], pc46[22], g45[22], ps45[22], pc45[22]);
FA1A GS45_23(ps46[22], pc46[23], g45[23], ps45[23], pc45[23]);
FA1A GS45_24(ps46[23], pc46[24], g45[24], ps45[24], pc45[24]);
FA1A GS45_25(ps46[24], pc46[25], g45[25], ps45[25], pc45[25]);
FA1A GS45_26(ps46[25], pc46[26], g45[26], ps45[26], pc45[26]);
FA1A GS45_27(ps46[26], pc46[27], g45[27], ps45[27], pc45[27]);
FA1A GS45_28(ps46[27], pc46[28], g45[28], ps45[28], pc45[28]);
FA1A GS45_29(ps46[28], pc46[29], g45[29], ps45[29], pc45[29]);
FA1A GS45_30(ps46[29], pc46[30], g45[30], ps45[30], pc45[30]);
FA1A GS45_31(ps46[30], pc46[31], g45[31], ps45[31], pc45[31]);
FA1A GS45_32(ps46[31], pc46[32], g45[32], ps45[32], pc45[32]);
FA1A GS45_33(ps46[32], pc46[33], g45[33], ps45[33], pc45[33]);
FA1A GS45_34(ps46[33], pc46[34], g45[34], ps45[34], pc45[34]);
FA1A GS45_35(ps46[34], pc46[35], g45[35], ps45[35], pc45[35]);
FA1A GS45_36(ps46[35], pc46[36], g45[36], ps45[36], pc45[36]);
FA1A GS45_37(ps46[36], pc46[37], g45[37], ps45[37], pc45[37]);
FA1A GS45_38(ps46[37], pc46[38], g45[38], ps45[38], pc45[38]);
FA1A GS45_39(ps46[38], pc46[39], g45[39], ps45[39], pc45[39]);
FA1A GS45_40(ps46[39], pc46[40], g45[40], ps45[40], pc45[40]);
FA1A GS45_41(ps46[40], pc46[41], g45[41], ps45[41], pc45[41]);
FA1A GS45_42(ps46[41], pc46[42], g45[42], ps45[42], pc45[42]);
FA1A GS45_43(ps46[42], pc46[43], g45[43], ps45[43], pc45[43]);
FA1A GS45_44(ps46[43], pc46[44], g45[44], ps45[44], pc45[44]);
FA1A GS45_45(ps46[44], pc46[45], g45[45], ps45[45], pc45[45]);
FA1A GS45_46(ps46[45], pc46[46], g45[46], ps45[46], pc45[46]);
FA1A GS45_47(ps46[46], pc46[47], g45[47], ps45[47], pc45[47]);
FA1A GS45_48(ps46[47], pc46[48], g45[48], ps45[48], pc45[48]);
FA1A GS45_49(ps46[48], pc46[49], g45[49], ps45[49], pc45[49]);
FA1A GS45_50(ps46[49], pc46[50], g45[50], ps45[50], pc45[50]);
FA1A GS45_51(ps46[50], pc46[51], g45[51], ps45[51], pc45[51]);
FA1A GS45_52(ps46[51], pc46[52], g45[52], ps45[52], pc45[52]);
FA1A GS45_53(ps46[52], pc46[53], g45[53], ps45[53], pc45[53]);
FA1A GS45_54(ps46[53], pc46[54], g45[54], ps45[54], pc45[54]);
FA1A GS45_55(ps46[54], pc46[55], g45[55], ps45[55], pc45[55]);
FA1A GS45_56(ps46[55], pc46[56], g45[56], ps45[56], pc45[56]);
FA1A GS45_57(ps46[56], pc46[57], g45[57], ps45[57], pc45[57]);
FA1A GS45_58(ps46[57], pc46[58], g45[58], ps45[58], pc45[58]);
FA1A GS45_59(ps46[58], pc46[59], g45[59], ps45[59], pc45[59]);
FA1A GS45_60(ps46[59], pc46[60], g45[60], ps45[60], pc45[60]);
FA1A GS45_61(ps46[60], pc46[61], g45[61], ps45[61], pc45[61]);
FA1A GS45_62(ps46[61], pc46[62], g45[62], ps45[62], pc45[62]);
FA1A GS45_63(ps46[62], pc46[63], g45[63], ps45[63], pc45[63]);
FA1A GS44_9(g45[8], pc45[9], g44[9], ps44[9], pc44[9]);
FA1A GS44_10(ps45[9], pc45[10], g44[10], ps44[10], pc44[10]);
FA1A GS44_11(ps45[10], pc45[11], g44[11], ps44[11], pc44[11]);
FA1A GS44_12(ps45[11], pc45[12], g44[12], ps44[12], pc44[12]);
FA1A GS44_13(ps45[12], pc45[13], g44[13], ps44[13], pc44[13]);
FA1A GS44_14(ps45[13], pc45[14], g44[14], ps44[14], pc44[14]);
FA1A GS44_15(ps45[14], pc45[15], g44[15], ps44[15], pc44[15]);
FA1A GS44_16(ps45[15], pc45[16], g44[16], ps44[16], pc44[16]);
FA1A GS44_17(ps45[16], pc45[17], g44[17], ps44[17], pc44[17]);
FA1A GS44_18(ps45[17], pc45[18], g44[18], ps44[18], pc44[18]);
FA1A GS44_19(ps45[18], pc45[19], g44[19], ps44[19], pc44[19]);
FA1A GS44_20(ps45[19], pc45[20], g44[20], ps44[20], pc44[20]);
FA1A GS44_21(ps45[20], pc45[21], g44[21], ps44[21], pc44[21]);
FA1A GS44_22(ps45[21], pc45[22], g44[22], ps44[22], pc44[22]);
FA1A GS44_23(ps45[22], pc45[23], g44[23], ps44[23], pc44[23]);
FA1A GS44_24(ps45[23], pc45[24], g44[24], ps44[24], pc44[24]);
FA1A GS44_25(ps45[24], pc45[25], g44[25], ps44[25], pc44[25]);
FA1A GS44_26(ps45[25], pc45[26], g44[26], ps44[26], pc44[26]);
FA1A GS44_27(ps45[26], pc45[27], g44[27], ps44[27], pc44[27]);
FA1A GS44_28(ps45[27], pc45[28], g44[28], ps44[28], pc44[28]);
FA1A GS44_29(ps45[28], pc45[29], g44[29], ps44[29], pc44[29]);
FA1A GS44_30(ps45[29], pc45[30], g44[30], ps44[30], pc44[30]);
FA1A GS44_31(ps45[30], pc45[31], g44[31], ps44[31], pc44[31]);
FA1A GS44_32(ps45[31], pc45[32], g44[32], ps44[32], pc44[32]);
FA1A GS44_33(ps45[32], pc45[33], g44[33], ps44[33], pc44[33]);
FA1A GS44_34(ps45[33], pc45[34], g44[34], ps44[34], pc44[34]);
FA1A GS44_35(ps45[34], pc45[35], g44[35], ps44[35], pc44[35]);
FA1A GS44_36(ps45[35], pc45[36], g44[36], ps44[36], pc44[36]);
FA1A GS44_37(ps45[36], pc45[37], g44[37], ps44[37], pc44[37]);
FA1A GS44_38(ps45[37], pc45[38], g44[38], ps44[38], pc44[38]);
FA1A GS44_39(ps45[38], pc45[39], g44[39], ps44[39], pc44[39]);
FA1A GS44_40(ps45[39], pc45[40], g44[40], ps44[40], pc44[40]);
FA1A GS44_41(ps45[40], pc45[41], g44[41], ps44[41], pc44[41]);
FA1A GS44_42(ps45[41], pc45[42], g44[42], ps44[42], pc44[42]);
FA1A GS44_43(ps45[42], pc45[43], g44[43], ps44[43], pc44[43]);
FA1A GS44_44(ps45[43], pc45[44], g44[44], ps44[44], pc44[44]);
FA1A GS44_45(ps45[44], pc45[45], g44[45], ps44[45], pc44[45]);
FA1A GS44_46(ps45[45], pc45[46], g44[46], ps44[46], pc44[46]);
FA1A GS44_47(ps45[46], pc45[47], g44[47], ps44[47], pc44[47]);
FA1A GS44_48(ps45[47], pc45[48], g44[48], ps44[48], pc44[48]);
FA1A GS44_49(ps45[48], pc45[49], g44[49], ps44[49], pc44[49]);
FA1A GS44_50(ps45[49], pc45[50], g44[50], ps44[50], pc44[50]);
FA1A GS44_51(ps45[50], pc45[51], g44[51], ps44[51], pc44[51]);
FA1A GS44_52(ps45[51], pc45[52], g44[52], ps44[52], pc44[52]);
FA1A GS44_53(ps45[52], pc45[53], g44[53], ps44[53], pc44[53]);
FA1A GS44_54(ps45[53], pc45[54], g44[54], ps44[54], pc44[54]);
FA1A GS44_55(ps45[54], pc45[55], g44[55], ps44[55], pc44[55]);
FA1A GS44_56(ps45[55], pc45[56], g44[56], ps44[56], pc44[56]);
FA1A GS44_57(ps45[56], pc45[57], g44[57], ps44[57], pc44[57]);
FA1A GS44_58(ps45[57], pc45[58], g44[58], ps44[58], pc44[58]);
FA1A GS44_59(ps45[58], pc45[59], g44[59], ps44[59], pc44[59]);
FA1A GS44_60(ps45[59], pc45[60], g44[60], ps44[60], pc44[60]);
FA1A GS44_61(ps45[60], pc45[61], g44[61], ps44[61], pc44[61]);
FA1A GS44_62(ps45[61], pc45[62], g44[62], ps44[62], pc44[62]);
FA1A GS44_63(ps45[62], pc45[63], g44[63], ps44[63], pc44[63]);
FA1A GS43_9(g44[8], pc44[9], g43[9], ps43[9], pc43[9]);
FA1A GS43_10(ps44[9], pc44[10], g43[10], ps43[10], pc43[10]);
FA1A GS43_11(ps44[10], pc44[11], g43[11], ps43[11], pc43[11]);
FA1A GS43_12(ps44[11], pc44[12], g43[12], ps43[12], pc43[12]);
FA1A GS43_13(ps44[12], pc44[13], g43[13], ps43[13], pc43[13]);
FA1A GS43_14(ps44[13], pc44[14], g43[14], ps43[14], pc43[14]);
FA1A GS43_15(ps44[14], pc44[15], g43[15], ps43[15], pc43[15]);
FA1A GS43_16(ps44[15], pc44[16], g43[16], ps43[16], pc43[16]);
FA1A GS43_17(ps44[16], pc44[17], g43[17], ps43[17], pc43[17]);
FA1A GS43_18(ps44[17], pc44[18], g43[18], ps43[18], pc43[18]);
FA1A GS43_19(ps44[18], pc44[19], g43[19], ps43[19], pc43[19]);
FA1A GS43_20(ps44[19], pc44[20], g43[20], ps43[20], pc43[20]);
FA1A GS43_21(ps44[20], pc44[21], g43[21], ps43[21], pc43[21]);
FA1A GS43_22(ps44[21], pc44[22], g43[22], ps43[22], pc43[22]);
FA1A GS43_23(ps44[22], pc44[23], g43[23], ps43[23], pc43[23]);
FA1A GS43_24(ps44[23], pc44[24], g43[24], ps43[24], pc43[24]);
FA1A GS43_25(ps44[24], pc44[25], g43[25], ps43[25], pc43[25]);
FA1A GS43_26(ps44[25], pc44[26], g43[26], ps43[26], pc43[26]);
FA1A GS43_27(ps44[26], pc44[27], g43[27], ps43[27], pc43[27]);
FA1A GS43_28(ps44[27], pc44[28], g43[28], ps43[28], pc43[28]);
FA1A GS43_29(ps44[28], pc44[29], g43[29], ps43[29], pc43[29]);
FA1A GS43_30(ps44[29], pc44[30], g43[30], ps43[30], pc43[30]);
FA1A GS43_31(ps44[30], pc44[31], g43[31], ps43[31], pc43[31]);
FA1A GS43_32(ps44[31], pc44[32], g43[32], ps43[32], pc43[32]);
FA1A GS43_33(ps44[32], pc44[33], g43[33], ps43[33], pc43[33]);
FA1A GS43_34(ps44[33], pc44[34], g43[34], ps43[34], pc43[34]);
FA1A GS43_35(ps44[34], pc44[35], g43[35], ps43[35], pc43[35]);
FA1A GS43_36(ps44[35], pc44[36], g43[36], ps43[36], pc43[36]);
FA1A GS43_37(ps44[36], pc44[37], g43[37], ps43[37], pc43[37]);
FA1A GS43_38(ps44[37], pc44[38], g43[38], ps43[38], pc43[38]);
FA1A GS43_39(ps44[38], pc44[39], g43[39], ps43[39], pc43[39]);
FA1A GS43_40(ps44[39], pc44[40], g43[40], ps43[40], pc43[40]);
FA1A GS43_41(ps44[40], pc44[41], g43[41], ps43[41], pc43[41]);
FA1A GS43_42(ps44[41], pc44[42], g43[42], ps43[42], pc43[42]);
FA1A GS43_43(ps44[42], pc44[43], g43[43], ps43[43], pc43[43]);
FA1A GS43_44(ps44[43], pc44[44], g43[44], ps43[44], pc43[44]);
FA1A GS43_45(ps44[44], pc44[45], g43[45], ps43[45], pc43[45]);
FA1A GS43_46(ps44[45], pc44[46], g43[46], ps43[46], pc43[46]);
FA1A GS43_47(ps44[46], pc44[47], g43[47], ps43[47], pc43[47]);
FA1A GS43_48(ps44[47], pc44[48], g43[48], ps43[48], pc43[48]);
FA1A GS43_49(ps44[48], pc44[49], g43[49], ps43[49], pc43[49]);
FA1A GS43_50(ps44[49], pc44[50], g43[50], ps43[50], pc43[50]);
FA1A GS43_51(ps44[50], pc44[51], g43[51], ps43[51], pc43[51]);
FA1A GS43_52(ps44[51], pc44[52], g43[52], ps43[52], pc43[52]);
FA1A GS43_53(ps44[52], pc44[53], g43[53], ps43[53], pc43[53]);
FA1A GS43_54(ps44[53], pc44[54], g43[54], ps43[54], pc43[54]);
FA1A GS43_55(ps44[54], pc44[55], g43[55], ps43[55], pc43[55]);
FA1A GS43_56(ps44[55], pc44[56], g43[56], ps43[56], pc43[56]);
FA1A GS43_57(ps44[56], pc44[57], g43[57], ps43[57], pc43[57]);
FA1A GS43_58(ps44[57], pc44[58], g43[58], ps43[58], pc43[58]);
FA1A GS43_59(ps44[58], pc44[59], g43[59], ps43[59], pc43[59]);
FA1A GS43_60(ps44[59], pc44[60], g43[60], ps43[60], pc43[60]);
FA1A GS43_61(ps44[60], pc44[61], g43[61], ps43[61], pc43[61]);
FA1A GS43_62(ps44[61], pc44[62], g43[62], ps43[62], pc43[62]);
FA1A GS43_63(ps44[62], pc44[63], g43[63], ps43[63], pc43[63]);
FA1A GS42_9(g43[8], pc43[9], g42[9], ps42[9], pc42[9]);
FA1A GS42_10(ps43[9], pc43[10], g42[10], ps42[10], pc42[10]);
FA1A GS42_11(ps43[10], pc43[11], g42[11], ps42[11], pc42[11]);
FA1A GS42_12(ps43[11], pc43[12], g42[12], ps42[12], pc42[12]);
FA1A GS42_13(ps43[12], pc43[13], g42[13], ps42[13], pc42[13]);
FA1A GS42_14(ps43[13], pc43[14], g42[14], ps42[14], pc42[14]);
FA1A GS42_15(ps43[14], pc43[15], g42[15], ps42[15], pc42[15]);
FA1A GS42_16(ps43[15], pc43[16], g42[16], ps42[16], pc42[16]);
FA1A GS42_17(ps43[16], pc43[17], g42[17], ps42[17], pc42[17]);
FA1A GS42_18(ps43[17], pc43[18], g42[18], ps42[18], pc42[18]);
FA1A GS42_19(ps43[18], pc43[19], g42[19], ps42[19], pc42[19]);
FA1A GS42_20(ps43[19], pc43[20], g42[20], ps42[20], pc42[20]);
FA1A GS42_21(ps43[20], pc43[21], g42[21], ps42[21], pc42[21]);
FA1A GS42_22(ps43[21], pc43[22], g42[22], ps42[22], pc42[22]);
FA1A GS42_23(ps43[22], pc43[23], g42[23], ps42[23], pc42[23]);
FA1A GS42_24(ps43[23], pc43[24], g42[24], ps42[24], pc42[24]);
FA1A GS42_25(ps43[24], pc43[25], g42[25], ps42[25], pc42[25]);
FA1A GS42_26(ps43[25], pc43[26], g42[26], ps42[26], pc42[26]);
FA1A GS42_27(ps43[26], pc43[27], g42[27], ps42[27], pc42[27]);
FA1A GS42_28(ps43[27], pc43[28], g42[28], ps42[28], pc42[28]);
FA1A GS42_29(ps43[28], pc43[29], g42[29], ps42[29], pc42[29]);
FA1A GS42_30(ps43[29], pc43[30], g42[30], ps42[30], pc42[30]);
FA1A GS42_31(ps43[30], pc43[31], g42[31], ps42[31], pc42[31]);
FA1A GS42_32(ps43[31], pc43[32], g42[32], ps42[32], pc42[32]);
FA1A GS42_33(ps43[32], pc43[33], g42[33], ps42[33], pc42[33]);
FA1A GS42_34(ps43[33], pc43[34], g42[34], ps42[34], pc42[34]);
FA1A GS42_35(ps43[34], pc43[35], g42[35], ps42[35], pc42[35]);
FA1A GS42_36(ps43[35], pc43[36], g42[36], ps42[36], pc42[36]);
FA1A GS42_37(ps43[36], pc43[37], g42[37], ps42[37], pc42[37]);
FA1A GS42_38(ps43[37], pc43[38], g42[38], ps42[38], pc42[38]);
FA1A GS42_39(ps43[38], pc43[39], g42[39], ps42[39], pc42[39]);
FA1A GS42_40(ps43[39], pc43[40], g42[40], ps42[40], pc42[40]);
FA1A GS42_41(ps43[40], pc43[41], g42[41], ps42[41], pc42[41]);
FA1A GS42_42(ps43[41], pc43[42], g42[42], ps42[42], pc42[42]);
FA1A GS42_43(ps43[42], pc43[43], g42[43], ps42[43], pc42[43]);
FA1A GS42_44(ps43[43], pc43[44], g42[44], ps42[44], pc42[44]);
FA1A GS42_45(ps43[44], pc43[45], g42[45], ps42[45], pc42[45]);
FA1A GS42_46(ps43[45], pc43[46], g42[46], ps42[46], pc42[46]);
FA1A GS42_47(ps43[46], pc43[47], g42[47], ps42[47], pc42[47]);
FA1A GS42_48(ps43[47], pc43[48], g42[48], ps42[48], pc42[48]);
FA1A GS42_49(ps43[48], pc43[49], g42[49], ps42[49], pc42[49]);
FA1A GS42_50(ps43[49], pc43[50], g42[50], ps42[50], pc42[50]);
FA1A GS42_51(ps43[50], pc43[51], g42[51], ps42[51], pc42[51]);
FA1A GS42_52(ps43[51], pc43[52], g42[52], ps42[52], pc42[52]);
FA1A GS42_53(ps43[52], pc43[53], g42[53], ps42[53], pc42[53]);
FA1A GS42_54(ps43[53], pc43[54], g42[54], ps42[54], pc42[54]);
FA1A GS42_55(ps43[54], pc43[55], g42[55], ps42[55], pc42[55]);
FA1A GS42_56(ps43[55], pc43[56], g42[56], ps42[56], pc42[56]);
FA1A GS42_57(ps43[56], pc43[57], g42[57], ps42[57], pc42[57]);
FA1A GS42_58(ps43[57], pc43[58], g42[58], ps42[58], pc42[58]);
FA1A GS42_59(ps43[58], pc43[59], g42[59], ps42[59], pc42[59]);
FA1A GS42_60(ps43[59], pc43[60], g42[60], ps42[60], pc42[60]);
FA1A GS42_61(ps43[60], pc43[61], g42[61], ps42[61], pc42[61]);
FA1A GS42_62(ps43[61], pc43[62], g42[62], ps42[62], pc42[62]);
FA1A GS42_63(ps43[62], pc43[63], g42[63], ps42[63], pc42[63]);
FA1A GS41_9(g42[8], pc42[9], g41[9], ps41[9], pc41[9]);
FA1A GS41_10(ps42[9], pc42[10], g41[10], ps41[10], pc41[10]);
FA1A GS41_11(ps42[10], pc42[11], g41[11], ps41[11], pc41[11]);
FA1A GS41_12(ps42[11], pc42[12], g41[12], ps41[12], pc41[12]);
FA1A GS41_13(ps42[12], pc42[13], g41[13], ps41[13], pc41[13]);
FA1A GS41_14(ps42[13], pc42[14], g41[14], ps41[14], pc41[14]);
FA1A GS41_15(ps42[14], pc42[15], g41[15], ps41[15], pc41[15]);
FA1A GS41_16(ps42[15], pc42[16], g41[16], ps41[16], pc41[16]);
FA1A GS41_17(ps42[16], pc42[17], g41[17], ps41[17], pc41[17]);
FA1A GS41_18(ps42[17], pc42[18], g41[18], ps41[18], pc41[18]);
FA1A GS41_19(ps42[18], pc42[19], g41[19], ps41[19], pc41[19]);
FA1A GS41_20(ps42[19], pc42[20], g41[20], ps41[20], pc41[20]);
FA1A GS41_21(ps42[20], pc42[21], g41[21], ps41[21], pc41[21]);
FA1A GS41_22(ps42[21], pc42[22], g41[22], ps41[22], pc41[22]);
FA1A GS41_23(ps42[22], pc42[23], g41[23], ps41[23], pc41[23]);
FA1A GS41_24(ps42[23], pc42[24], g41[24], ps41[24], pc41[24]);
FA1A GS41_25(ps42[24], pc42[25], g41[25], ps41[25], pc41[25]);
FA1A GS41_26(ps42[25], pc42[26], g41[26], ps41[26], pc41[26]);
FA1A GS41_27(ps42[26], pc42[27], g41[27], ps41[27], pc41[27]);
FA1A GS41_28(ps42[27], pc42[28], g41[28], ps41[28], pc41[28]);
FA1A GS41_29(ps42[28], pc42[29], g41[29], ps41[29], pc41[29]);
FA1A GS41_30(ps42[29], pc42[30], g41[30], ps41[30], pc41[30]);
FA1A GS41_31(ps42[30], pc42[31], g41[31], ps41[31], pc41[31]);
FA1A GS41_32(ps42[31], pc42[32], g41[32], ps41[32], pc41[32]);
FA1A GS41_33(ps42[32], pc42[33], g41[33], ps41[33], pc41[33]);
FA1A GS41_34(ps42[33], pc42[34], g41[34], ps41[34], pc41[34]);
FA1A GS41_35(ps42[34], pc42[35], g41[35], ps41[35], pc41[35]);
FA1A GS41_36(ps42[35], pc42[36], g41[36], ps41[36], pc41[36]);
FA1A GS41_37(ps42[36], pc42[37], g41[37], ps41[37], pc41[37]);
FA1A GS41_38(ps42[37], pc42[38], g41[38], ps41[38], pc41[38]);
FA1A GS41_39(ps42[38], pc42[39], g41[39], ps41[39], pc41[39]);
FA1A GS41_40(ps42[39], pc42[40], g41[40], ps41[40], pc41[40]);
FA1A GS41_41(ps42[40], pc42[41], g41[41], ps41[41], pc41[41]);
FA1A GS41_42(ps42[41], pc42[42], g41[42], ps41[42], pc41[42]);
FA1A GS41_43(ps42[42], pc42[43], g41[43], ps41[43], pc41[43]);
FA1A GS41_44(ps42[43], pc42[44], g41[44], ps41[44], pc41[44]);
FA1A GS41_45(ps42[44], pc42[45], g41[45], ps41[45], pc41[45]);
FA1A GS41_46(ps42[45], pc42[46], g41[46], ps41[46], pc41[46]);
FA1A GS41_47(ps42[46], pc42[47], g41[47], ps41[47], pc41[47]);
FA1A GS41_48(ps42[47], pc42[48], g41[48], ps41[48], pc41[48]);
FA1A GS41_49(ps42[48], pc42[49], g41[49], ps41[49], pc41[49]);
FA1A GS41_50(ps42[49], pc42[50], g41[50], ps41[50], pc41[50]);
FA1A GS41_51(ps42[50], pc42[51], g41[51], ps41[51], pc41[51]);
FA1A GS41_52(ps42[51], pc42[52], g41[52], ps41[52], pc41[52]);
FA1A GS41_53(ps42[52], pc42[53], g41[53], ps41[53], pc41[53]);
FA1A GS41_54(ps42[53], pc42[54], g41[54], ps41[54], pc41[54]);
FA1A GS41_55(ps42[54], pc42[55], g41[55], ps41[55], pc41[55]);
FA1A GS41_56(ps42[55], pc42[56], g41[56], ps41[56], pc41[56]);
FA1A GS41_57(ps42[56], pc42[57], g41[57], ps41[57], pc41[57]);
FA1A GS41_58(ps42[57], pc42[58], g41[58], ps41[58], pc41[58]);
FA1A GS41_59(ps42[58], pc42[59], g41[59], ps41[59], pc41[59]);
FA1A GS41_60(ps42[59], pc42[60], g41[60], ps41[60], pc41[60]);
FA1A GS41_61(ps42[60], pc42[61], g41[61], ps41[61], pc41[61]);
FA1A GS41_62(ps42[61], pc42[62], g41[62], ps41[62], pc41[62]);
FA1A GS41_63(ps42[62], pc42[63], g41[63], ps41[63], pc41[63]);
FA1A GS40_9(g41[8], pc41[9], g40[9], ps40[9], pc40[9]);
FA1A GS40_10(ps41[9], pc41[10], g40[10], ps40[10], pc40[10]);
FA1A GS40_11(ps41[10], pc41[11], g40[11], ps40[11], pc40[11]);
FA1A GS40_12(ps41[11], pc41[12], g40[12], ps40[12], pc40[12]);
FA1A GS40_13(ps41[12], pc41[13], g40[13], ps40[13], pc40[13]);
FA1A GS40_14(ps41[13], pc41[14], g40[14], ps40[14], pc40[14]);
FA1A GS40_15(ps41[14], pc41[15], g40[15], ps40[15], pc40[15]);
FA1A GS40_16(ps41[15], pc41[16], g40[16], ps40[16], pc40[16]);
FA1A GS40_17(ps41[16], pc41[17], g40[17], ps40[17], pc40[17]);
FA1A GS40_18(ps41[17], pc41[18], g40[18], ps40[18], pc40[18]);
FA1A GS40_19(ps41[18], pc41[19], g40[19], ps40[19], pc40[19]);
FA1A GS40_20(ps41[19], pc41[20], g40[20], ps40[20], pc40[20]);
FA1A GS40_21(ps41[20], pc41[21], g40[21], ps40[21], pc40[21]);
FA1A GS40_22(ps41[21], pc41[22], g40[22], ps40[22], pc40[22]);
FA1A GS40_23(ps41[22], pc41[23], g40[23], ps40[23], pc40[23]);
FA1A GS40_24(ps41[23], pc41[24], g40[24], ps40[24], pc40[24]);
FA1A GS40_25(ps41[24], pc41[25], g40[25], ps40[25], pc40[25]);
FA1A GS40_26(ps41[25], pc41[26], g40[26], ps40[26], pc40[26]);
FA1A GS40_27(ps41[26], pc41[27], g40[27], ps40[27], pc40[27]);
FA1A GS40_28(ps41[27], pc41[28], g40[28], ps40[28], pc40[28]);
FA1A GS40_29(ps41[28], pc41[29], g40[29], ps40[29], pc40[29]);
FA1A GS40_30(ps41[29], pc41[30], g40[30], ps40[30], pc40[30]);
FA1A GS40_31(ps41[30], pc41[31], g40[31], ps40[31], pc40[31]);
FA1A GS40_32(ps41[31], pc41[32], g40[32], ps40[32], pc40[32]);
FA1A GS40_33(ps41[32], pc41[33], g40[33], ps40[33], pc40[33]);
FA1A GS40_34(ps41[33], pc41[34], g40[34], ps40[34], pc40[34]);
FA1A GS40_35(ps41[34], pc41[35], g40[35], ps40[35], pc40[35]);
FA1A GS40_36(ps41[35], pc41[36], g40[36], ps40[36], pc40[36]);
FA1A GS40_37(ps41[36], pc41[37], g40[37], ps40[37], pc40[37]);
FA1A GS40_38(ps41[37], pc41[38], g40[38], ps40[38], pc40[38]);
FA1A GS40_39(ps41[38], pc41[39], g40[39], ps40[39], pc40[39]);
FA1A GS40_40(ps41[39], pc41[40], g40[40], ps40[40], pc40[40]);
FA1A GS40_41(ps41[40], pc41[41], g40[41], ps40[41], pc40[41]);
FA1A GS40_42(ps41[41], pc41[42], g40[42], ps40[42], pc40[42]);
FA1A GS40_43(ps41[42], pc41[43], g40[43], ps40[43], pc40[43]);
FA1A GS40_44(ps41[43], pc41[44], g40[44], ps40[44], pc40[44]);
FA1A GS40_45(ps41[44], pc41[45], g40[45], ps40[45], pc40[45]);
FA1A GS40_46(ps41[45], pc41[46], g40[46], ps40[46], pc40[46]);
FA1A GS40_47(ps41[46], pc41[47], g40[47], ps40[47], pc40[47]);
FA1A GS40_48(ps41[47], pc41[48], g40[48], ps40[48], pc40[48]);
FA1A GS40_49(ps41[48], pc41[49], g40[49], ps40[49], pc40[49]);
FA1A GS40_50(ps41[49], pc41[50], g40[50], ps40[50], pc40[50]);
FA1A GS40_51(ps41[50], pc41[51], g40[51], ps40[51], pc40[51]);
FA1A GS40_52(ps41[51], pc41[52], g40[52], ps40[52], pc40[52]);
FA1A GS40_53(ps41[52], pc41[53], g40[53], ps40[53], pc40[53]);
FA1A GS40_54(ps41[53], pc41[54], g40[54], ps40[54], pc40[54]);
FA1A GS40_55(ps41[54], pc41[55], g40[55], ps40[55], pc40[55]);
FA1A GS40_56(ps41[55], pc41[56], g40[56], ps40[56], pc40[56]);
FA1A GS40_57(ps41[56], pc41[57], g40[57], ps40[57], pc40[57]);
FA1A GS40_58(ps41[57], pc41[58], g40[58], ps40[58], pc40[58]);
FA1A GS40_59(ps41[58], pc41[59], g40[59], ps40[59], pc40[59]);
FA1A GS40_60(ps41[59], pc41[60], g40[60], ps40[60], pc40[60]);
FA1A GS40_61(ps41[60], pc41[61], g40[61], ps40[61], pc40[61]);
FA1A GS40_62(ps41[61], pc41[62], g40[62], ps40[62], pc40[62]);
FA1A GS40_63(ps41[62], pc41[63], g40[63], ps40[63], pc40[63]);
FA1A GS39_9(g40[8], pc40[9], g39[9], ps39[9], pc39[9]);
FA1A GS39_10(ps40[9], pc40[10], g39[10], ps39[10], pc39[10]);
FA1A GS39_11(ps40[10], pc40[11], g39[11], ps39[11], pc39[11]);
FA1A GS39_12(ps40[11], pc40[12], g39[12], ps39[12], pc39[12]);
FA1A GS39_13(ps40[12], pc40[13], g39[13], ps39[13], pc39[13]);
FA1A GS39_14(ps40[13], pc40[14], g39[14], ps39[14], pc39[14]);
FA1A GS39_15(ps40[14], pc40[15], g39[15], ps39[15], pc39[15]);
FA1A GS39_16(ps40[15], pc40[16], g39[16], ps39[16], pc39[16]);
FA1A GS39_17(ps40[16], pc40[17], g39[17], ps39[17], pc39[17]);
FA1A GS39_18(ps40[17], pc40[18], g39[18], ps39[18], pc39[18]);
FA1A GS39_19(ps40[18], pc40[19], g39[19], ps39[19], pc39[19]);
FA1A GS39_20(ps40[19], pc40[20], g39[20], ps39[20], pc39[20]);
FA1A GS39_21(ps40[20], pc40[21], g39[21], ps39[21], pc39[21]);
FA1A GS39_22(ps40[21], pc40[22], g39[22], ps39[22], pc39[22]);
FA1A GS39_23(ps40[22], pc40[23], g39[23], ps39[23], pc39[23]);
FA1A GS39_24(ps40[23], pc40[24], g39[24], ps39[24], pc39[24]);
FA1A GS39_25(ps40[24], pc40[25], g39[25], ps39[25], pc39[25]);
FA1A GS39_26(ps40[25], pc40[26], g39[26], ps39[26], pc39[26]);
FA1A GS39_27(ps40[26], pc40[27], g39[27], ps39[27], pc39[27]);
FA1A GS39_28(ps40[27], pc40[28], g39[28], ps39[28], pc39[28]);
FA1A GS39_29(ps40[28], pc40[29], g39[29], ps39[29], pc39[29]);
FA1A GS39_30(ps40[29], pc40[30], g39[30], ps39[30], pc39[30]);
FA1A GS39_31(ps40[30], pc40[31], g39[31], ps39[31], pc39[31]);
FA1A GS39_32(ps40[31], pc40[32], g39[32], ps39[32], pc39[32]);
FA1A GS39_33(ps40[32], pc40[33], g39[33], ps39[33], pc39[33]);
FA1A GS39_34(ps40[33], pc40[34], g39[34], ps39[34], pc39[34]);
FA1A GS39_35(ps40[34], pc40[35], g39[35], ps39[35], pc39[35]);
FA1A GS39_36(ps40[35], pc40[36], g39[36], ps39[36], pc39[36]);
FA1A GS39_37(ps40[36], pc40[37], g39[37], ps39[37], pc39[37]);
FA1A GS39_38(ps40[37], pc40[38], g39[38], ps39[38], pc39[38]);
FA1A GS39_39(ps40[38], pc40[39], g39[39], ps39[39], pc39[39]);
FA1A GS39_40(ps40[39], pc40[40], g39[40], ps39[40], pc39[40]);
FA1A GS39_41(ps40[40], pc40[41], g39[41], ps39[41], pc39[41]);
FA1A GS39_42(ps40[41], pc40[42], g39[42], ps39[42], pc39[42]);
FA1A GS39_43(ps40[42], pc40[43], g39[43], ps39[43], pc39[43]);
FA1A GS39_44(ps40[43], pc40[44], g39[44], ps39[44], pc39[44]);
FA1A GS39_45(ps40[44], pc40[45], g39[45], ps39[45], pc39[45]);
FA1A GS39_46(ps40[45], pc40[46], g39[46], ps39[46], pc39[46]);
FA1A GS39_47(ps40[46], pc40[47], g39[47], ps39[47], pc39[47]);
FA1A GS39_48(ps40[47], pc40[48], g39[48], ps39[48], pc39[48]);
FA1A GS39_49(ps40[48], pc40[49], g39[49], ps39[49], pc39[49]);
FA1A GS39_50(ps40[49], pc40[50], g39[50], ps39[50], pc39[50]);
FA1A GS39_51(ps40[50], pc40[51], g39[51], ps39[51], pc39[51]);
FA1A GS39_52(ps40[51], pc40[52], g39[52], ps39[52], pc39[52]);
FA1A GS39_53(ps40[52], pc40[53], g39[53], ps39[53], pc39[53]);
FA1A GS39_54(ps40[53], pc40[54], g39[54], ps39[54], pc39[54]);
FA1A GS39_55(ps40[54], pc40[55], g39[55], ps39[55], pc39[55]);
FA1A GS39_56(ps40[55], pc40[56], g39[56], ps39[56], pc39[56]);
FA1A GS39_57(ps40[56], pc40[57], g39[57], ps39[57], pc39[57]);
FA1A GS39_58(ps40[57], pc40[58], g39[58], ps39[58], pc39[58]);
FA1A GS39_59(ps40[58], pc40[59], g39[59], ps39[59], pc39[59]);
FA1A GS39_60(ps40[59], pc40[60], g39[60], ps39[60], pc39[60]);
FA1A GS39_61(ps40[60], pc40[61], g39[61], ps39[61], pc39[61]);
FA1A GS39_62(ps40[61], pc40[62], g39[62], ps39[62], pc39[62]);
FA1A GS39_63(ps40[62], pc40[63], g39[63], ps39[63], pc39[63]);
FA1A GS38_9(g39[8], pc39[9], g38[9], ps38[9], pc38[9]);
FA1A GS38_10(ps39[9], pc39[10], g38[10], ps38[10], pc38[10]);
FA1A GS38_11(ps39[10], pc39[11], g38[11], ps38[11], pc38[11]);
FA1A GS38_12(ps39[11], pc39[12], g38[12], ps38[12], pc38[12]);
FA1A GS38_13(ps39[12], pc39[13], g38[13], ps38[13], pc38[13]);
FA1A GS38_14(ps39[13], pc39[14], g38[14], ps38[14], pc38[14]);
FA1A GS38_15(ps39[14], pc39[15], g38[15], ps38[15], pc38[15]);
FA1A GS38_16(ps39[15], pc39[16], g38[16], ps38[16], pc38[16]);
FA1A GS38_17(ps39[16], pc39[17], g38[17], ps38[17], pc38[17]);
FA1A GS38_18(ps39[17], pc39[18], g38[18], ps38[18], pc38[18]);
FA1A GS38_19(ps39[18], pc39[19], g38[19], ps38[19], pc38[19]);
FA1A GS38_20(ps39[19], pc39[20], g38[20], ps38[20], pc38[20]);
FA1A GS38_21(ps39[20], pc39[21], g38[21], ps38[21], pc38[21]);
FA1A GS38_22(ps39[21], pc39[22], g38[22], ps38[22], pc38[22]);
FA1A GS38_23(ps39[22], pc39[23], g38[23], ps38[23], pc38[23]);
FA1A GS38_24(ps39[23], pc39[24], g38[24], ps38[24], pc38[24]);
FA1A GS38_25(ps39[24], pc39[25], g38[25], ps38[25], pc38[25]);
FA1A GS38_26(ps39[25], pc39[26], g38[26], ps38[26], pc38[26]);
FA1A GS38_27(ps39[26], pc39[27], g38[27], ps38[27], pc38[27]);
FA1A GS38_28(ps39[27], pc39[28], g38[28], ps38[28], pc38[28]);
FA1A GS38_29(ps39[28], pc39[29], g38[29], ps38[29], pc38[29]);
FA1A GS38_30(ps39[29], pc39[30], g38[30], ps38[30], pc38[30]);
FA1A GS38_31(ps39[30], pc39[31], g38[31], ps38[31], pc38[31]);
FA1A GS38_32(ps39[31], pc39[32], g38[32], ps38[32], pc38[32]);
FA1A GS38_33(ps39[32], pc39[33], g38[33], ps38[33], pc38[33]);
FA1A GS38_34(ps39[33], pc39[34], g38[34], ps38[34], pc38[34]);
FA1A GS38_35(ps39[34], pc39[35], g38[35], ps38[35], pc38[35]);
FA1A GS38_36(ps39[35], pc39[36], g38[36], ps38[36], pc38[36]);
FA1A GS38_37(ps39[36], pc39[37], g38[37], ps38[37], pc38[37]);
FA1A GS38_38(ps39[37], pc39[38], g38[38], ps38[38], pc38[38]);
FA1A GS38_39(ps39[38], pc39[39], g38[39], ps38[39], pc38[39]);
FA1A GS38_40(ps39[39], pc39[40], g38[40], ps38[40], pc38[40]);
FA1A GS38_41(ps39[40], pc39[41], g38[41], ps38[41], pc38[41]);
FA1A GS38_42(ps39[41], pc39[42], g38[42], ps38[42], pc38[42]);
FA1A GS38_43(ps39[42], pc39[43], g38[43], ps38[43], pc38[43]);
FA1A GS38_44(ps39[43], pc39[44], g38[44], ps38[44], pc38[44]);
FA1A GS38_45(ps39[44], pc39[45], g38[45], ps38[45], pc38[45]);
FA1A GS38_46(ps39[45], pc39[46], g38[46], ps38[46], pc38[46]);
FA1A GS38_47(ps39[46], pc39[47], g38[47], ps38[47], pc38[47]);
FA1A GS38_48(ps39[47], pc39[48], g38[48], ps38[48], pc38[48]);
FA1A GS38_49(ps39[48], pc39[49], g38[49], ps38[49], pc38[49]);
FA1A GS38_50(ps39[49], pc39[50], g38[50], ps38[50], pc38[50]);
FA1A GS38_51(ps39[50], pc39[51], g38[51], ps38[51], pc38[51]);
FA1A GS38_52(ps39[51], pc39[52], g38[52], ps38[52], pc38[52]);
FA1A GS38_53(ps39[52], pc39[53], g38[53], ps38[53], pc38[53]);
FA1A GS38_54(ps39[53], pc39[54], g38[54], ps38[54], pc38[54]);
FA1A GS38_55(ps39[54], pc39[55], g38[55], ps38[55], pc38[55]);
FA1A GS38_56(ps39[55], pc39[56], g38[56], ps38[56], pc38[56]);
FA1A GS38_57(ps39[56], pc39[57], g38[57], ps38[57], pc38[57]);
FA1A GS38_58(ps39[57], pc39[58], g38[58], ps38[58], pc38[58]);
FA1A GS38_59(ps39[58], pc39[59], g38[59], ps38[59], pc38[59]);
FA1A GS38_60(ps39[59], pc39[60], g38[60], ps38[60], pc38[60]);
FA1A GS38_61(ps39[60], pc39[61], g38[61], ps38[61], pc38[61]);
FA1A GS38_62(ps39[61], pc39[62], g38[62], ps38[62], pc38[62]);
FA1A GS38_63(ps39[62], pc39[63], g38[63], ps38[63], pc38[63]);
FA1A GS37_9(g38[8], pc38[9], g37[9], ps37[9], pc37[9]);
FA1A GS37_10(ps38[9], pc38[10], g37[10], ps37[10], pc37[10]);
FA1A GS37_11(ps38[10], pc38[11], g37[11], ps37[11], pc37[11]);
FA1A GS37_12(ps38[11], pc38[12], g37[12], ps37[12], pc37[12]);
FA1A GS37_13(ps38[12], pc38[13], g37[13], ps37[13], pc37[13]);
FA1A GS37_14(ps38[13], pc38[14], g37[14], ps37[14], pc37[14]);
FA1A GS37_15(ps38[14], pc38[15], g37[15], ps37[15], pc37[15]);
FA1A GS37_16(ps38[15], pc38[16], g37[16], ps37[16], pc37[16]);
FA1A GS37_17(ps38[16], pc38[17], g37[17], ps37[17], pc37[17]);
FA1A GS37_18(ps38[17], pc38[18], g37[18], ps37[18], pc37[18]);
FA1A GS37_19(ps38[18], pc38[19], g37[19], ps37[19], pc37[19]);
FA1A GS37_20(ps38[19], pc38[20], g37[20], ps37[20], pc37[20]);
FA1A GS37_21(ps38[20], pc38[21], g37[21], ps37[21], pc37[21]);
FA1A GS37_22(ps38[21], pc38[22], g37[22], ps37[22], pc37[22]);
FA1A GS37_23(ps38[22], pc38[23], g37[23], ps37[23], pc37[23]);
FA1A GS37_24(ps38[23], pc38[24], g37[24], ps37[24], pc37[24]);
FA1A GS37_25(ps38[24], pc38[25], g37[25], ps37[25], pc37[25]);
FA1A GS37_26(ps38[25], pc38[26], g37[26], ps37[26], pc37[26]);
FA1A GS37_27(ps38[26], pc38[27], g37[27], ps37[27], pc37[27]);
FA1A GS37_28(ps38[27], pc38[28], g37[28], ps37[28], pc37[28]);
FA1A GS37_29(ps38[28], pc38[29], g37[29], ps37[29], pc37[29]);
FA1A GS37_30(ps38[29], pc38[30], g37[30], ps37[30], pc37[30]);
FA1A GS37_31(ps38[30], pc38[31], g37[31], ps37[31], pc37[31]);
FA1A GS37_32(ps38[31], pc38[32], g37[32], ps37[32], pc37[32]);
FA1A GS37_33(ps38[32], pc38[33], g37[33], ps37[33], pc37[33]);
FA1A GS37_34(ps38[33], pc38[34], g37[34], ps37[34], pc37[34]);
FA1A GS37_35(ps38[34], pc38[35], g37[35], ps37[35], pc37[35]);
FA1A GS37_36(ps38[35], pc38[36], g37[36], ps37[36], pc37[36]);
FA1A GS37_37(ps38[36], pc38[37], g37[37], ps37[37], pc37[37]);
FA1A GS37_38(ps38[37], pc38[38], g37[38], ps37[38], pc37[38]);
FA1A GS37_39(ps38[38], pc38[39], g37[39], ps37[39], pc37[39]);
FA1A GS37_40(ps38[39], pc38[40], g37[40], ps37[40], pc37[40]);
FA1A GS37_41(ps38[40], pc38[41], g37[41], ps37[41], pc37[41]);
FA1A GS37_42(ps38[41], pc38[42], g37[42], ps37[42], pc37[42]);
FA1A GS37_43(ps38[42], pc38[43], g37[43], ps37[43], pc37[43]);
FA1A GS37_44(ps38[43], pc38[44], g37[44], ps37[44], pc37[44]);
FA1A GS37_45(ps38[44], pc38[45], g37[45], ps37[45], pc37[45]);
FA1A GS37_46(ps38[45], pc38[46], g37[46], ps37[46], pc37[46]);
FA1A GS37_47(ps38[46], pc38[47], g37[47], ps37[47], pc37[47]);
FA1A GS37_48(ps38[47], pc38[48], g37[48], ps37[48], pc37[48]);
FA1A GS37_49(ps38[48], pc38[49], g37[49], ps37[49], pc37[49]);
FA1A GS37_50(ps38[49], pc38[50], g37[50], ps37[50], pc37[50]);
FA1A GS37_51(ps38[50], pc38[51], g37[51], ps37[51], pc37[51]);
FA1A GS37_52(ps38[51], pc38[52], g37[52], ps37[52], pc37[52]);
FA1A GS37_53(ps38[52], pc38[53], g37[53], ps37[53], pc37[53]);
FA1A GS37_54(ps38[53], pc38[54], g37[54], ps37[54], pc37[54]);
FA1A GS37_55(ps38[54], pc38[55], g37[55], ps37[55], pc37[55]);
FA1A GS37_56(ps38[55], pc38[56], g37[56], ps37[56], pc37[56]);
FA1A GS37_57(ps38[56], pc38[57], g37[57], ps37[57], pc37[57]);
FA1A GS37_58(ps38[57], pc38[58], g37[58], ps37[58], pc37[58]);
FA1A GS37_59(ps38[58], pc38[59], g37[59], ps37[59], pc37[59]);
FA1A GS37_60(ps38[59], pc38[60], g37[60], ps37[60], pc37[60]);
FA1A GS37_61(ps38[60], pc38[61], g37[61], ps37[61], pc37[61]);
FA1A GS37_62(ps38[61], pc38[62], g37[62], ps37[62], pc37[62]);
FA1A GS37_63(ps38[62], pc38[63], g37[63], ps37[63], pc37[63]);
FA1A GS36_9(g37[8], pc37[9], g36[9], ps36[9], pc36[9]);
FA1A GS36_10(ps37[9], pc37[10], g36[10], ps36[10], pc36[10]);
FA1A GS36_11(ps37[10], pc37[11], g36[11], ps36[11], pc36[11]);
FA1A GS36_12(ps37[11], pc37[12], g36[12], ps36[12], pc36[12]);
FA1A GS36_13(ps37[12], pc37[13], g36[13], ps36[13], pc36[13]);
FA1A GS36_14(ps37[13], pc37[14], g36[14], ps36[14], pc36[14]);
FA1A GS36_15(ps37[14], pc37[15], g36[15], ps36[15], pc36[15]);
FA1A GS36_16(ps37[15], pc37[16], g36[16], ps36[16], pc36[16]);
FA1A GS36_17(ps37[16], pc37[17], g36[17], ps36[17], pc36[17]);
FA1A GS36_18(ps37[17], pc37[18], g36[18], ps36[18], pc36[18]);
FA1A GS36_19(ps37[18], pc37[19], g36[19], ps36[19], pc36[19]);
FA1A GS36_20(ps37[19], pc37[20], g36[20], ps36[20], pc36[20]);
FA1A GS36_21(ps37[20], pc37[21], g36[21], ps36[21], pc36[21]);
FA1A GS36_22(ps37[21], pc37[22], g36[22], ps36[22], pc36[22]);
FA1A GS36_23(ps37[22], pc37[23], g36[23], ps36[23], pc36[23]);
FA1A GS36_24(ps37[23], pc37[24], g36[24], ps36[24], pc36[24]);
FA1A GS36_25(ps37[24], pc37[25], g36[25], ps36[25], pc36[25]);
FA1A GS36_26(ps37[25], pc37[26], g36[26], ps36[26], pc36[26]);
FA1A GS36_27(ps37[26], pc37[27], g36[27], ps36[27], pc36[27]);
FA1A GS36_28(ps37[27], pc37[28], g36[28], ps36[28], pc36[28]);
FA1A GS36_29(ps37[28], pc37[29], g36[29], ps36[29], pc36[29]);
FA1A GS36_30(ps37[29], pc37[30], g36[30], ps36[30], pc36[30]);
FA1A GS36_31(ps37[30], pc37[31], g36[31], ps36[31], pc36[31]);
FA1A GS36_32(ps37[31], pc37[32], g36[32], ps36[32], pc36[32]);
FA1A GS36_33(ps37[32], pc37[33], g36[33], ps36[33], pc36[33]);
FA1A GS36_34(ps37[33], pc37[34], g36[34], ps36[34], pc36[34]);
FA1A GS36_35(ps37[34], pc37[35], g36[35], ps36[35], pc36[35]);
FA1A GS36_36(ps37[35], pc37[36], g36[36], ps36[36], pc36[36]);
FA1A GS36_37(ps37[36], pc37[37], g36[37], ps36[37], pc36[37]);
FA1A GS36_38(ps37[37], pc37[38], g36[38], ps36[38], pc36[38]);
FA1A GS36_39(ps37[38], pc37[39], g36[39], ps36[39], pc36[39]);
FA1A GS36_40(ps37[39], pc37[40], g36[40], ps36[40], pc36[40]);
FA1A GS36_41(ps37[40], pc37[41], g36[41], ps36[41], pc36[41]);
FA1A GS36_42(ps37[41], pc37[42], g36[42], ps36[42], pc36[42]);
FA1A GS36_43(ps37[42], pc37[43], g36[43], ps36[43], pc36[43]);
FA1A GS36_44(ps37[43], pc37[44], g36[44], ps36[44], pc36[44]);
FA1A GS36_45(ps37[44], pc37[45], g36[45], ps36[45], pc36[45]);
FA1A GS36_46(ps37[45], pc37[46], g36[46], ps36[46], pc36[46]);
FA1A GS36_47(ps37[46], pc37[47], g36[47], ps36[47], pc36[47]);
FA1A GS36_48(ps37[47], pc37[48], g36[48], ps36[48], pc36[48]);
FA1A GS36_49(ps37[48], pc37[49], g36[49], ps36[49], pc36[49]);
FA1A GS36_50(ps37[49], pc37[50], g36[50], ps36[50], pc36[50]);
FA1A GS36_51(ps37[50], pc37[51], g36[51], ps36[51], pc36[51]);
FA1A GS36_52(ps37[51], pc37[52], g36[52], ps36[52], pc36[52]);
FA1A GS36_53(ps37[52], pc37[53], g36[53], ps36[53], pc36[53]);
FA1A GS36_54(ps37[53], pc37[54], g36[54], ps36[54], pc36[54]);
FA1A GS36_55(ps37[54], pc37[55], g36[55], ps36[55], pc36[55]);
FA1A GS36_56(ps37[55], pc37[56], g36[56], ps36[56], pc36[56]);
FA1A GS36_57(ps37[56], pc37[57], g36[57], ps36[57], pc36[57]);
FA1A GS36_58(ps37[57], pc37[58], g36[58], ps36[58], pc36[58]);
FA1A GS36_59(ps37[58], pc37[59], g36[59], ps36[59], pc36[59]);
FA1A GS36_60(ps37[59], pc37[60], g36[60], ps36[60], pc36[60]);
FA1A GS36_61(ps37[60], pc37[61], g36[61], ps36[61], pc36[61]);
FA1A GS36_62(ps37[61], pc37[62], g36[62], ps36[62], pc36[62]);
FA1A GS36_63(ps37[62], pc37[63], g36[63], ps36[63], pc36[63]);
FA1A GS35_9(g36[8], pc36[9], g35[9], ps35[9], pc35[9]);
FA1A GS35_10(ps36[9], pc36[10], g35[10], ps35[10], pc35[10]);
FA1A GS35_11(ps36[10], pc36[11], g35[11], ps35[11], pc35[11]);
FA1A GS35_12(ps36[11], pc36[12], g35[12], ps35[12], pc35[12]);
FA1A GS35_13(ps36[12], pc36[13], g35[13], ps35[13], pc35[13]);
FA1A GS35_14(ps36[13], pc36[14], g35[14], ps35[14], pc35[14]);
FA1A GS35_15(ps36[14], pc36[15], g35[15], ps35[15], pc35[15]);
FA1A GS35_16(ps36[15], pc36[16], g35[16], ps35[16], pc35[16]);
FA1A GS35_17(ps36[16], pc36[17], g35[17], ps35[17], pc35[17]);
FA1A GS35_18(ps36[17], pc36[18], g35[18], ps35[18], pc35[18]);
FA1A GS35_19(ps36[18], pc36[19], g35[19], ps35[19], pc35[19]);
FA1A GS35_20(ps36[19], pc36[20], g35[20], ps35[20], pc35[20]);
FA1A GS35_21(ps36[20], pc36[21], g35[21], ps35[21], pc35[21]);
FA1A GS35_22(ps36[21], pc36[22], g35[22], ps35[22], pc35[22]);
FA1A GS35_23(ps36[22], pc36[23], g35[23], ps35[23], pc35[23]);
FA1A GS35_24(ps36[23], pc36[24], g35[24], ps35[24], pc35[24]);
FA1A GS35_25(ps36[24], pc36[25], g35[25], ps35[25], pc35[25]);
FA1A GS35_26(ps36[25], pc36[26], g35[26], ps35[26], pc35[26]);
FA1A GS35_27(ps36[26], pc36[27], g35[27], ps35[27], pc35[27]);
FA1A GS35_28(ps36[27], pc36[28], g35[28], ps35[28], pc35[28]);
FA1A GS35_29(ps36[28], pc36[29], g35[29], ps35[29], pc35[29]);
FA1A GS35_30(ps36[29], pc36[30], g35[30], ps35[30], pc35[30]);
FA1A GS35_31(ps36[30], pc36[31], g35[31], ps35[31], pc35[31]);
FA1A GS35_32(ps36[31], pc36[32], g35[32], ps35[32], pc35[32]);
FA1A GS35_33(ps36[32], pc36[33], g35[33], ps35[33], pc35[33]);
FA1A GS35_34(ps36[33], pc36[34], g35[34], ps35[34], pc35[34]);
FA1A GS35_35(ps36[34], pc36[35], g35[35], ps35[35], pc35[35]);
FA1A GS35_36(ps36[35], pc36[36], g35[36], ps35[36], pc35[36]);
FA1A GS35_37(ps36[36], pc36[37], g35[37], ps35[37], pc35[37]);
FA1A GS35_38(ps36[37], pc36[38], g35[38], ps35[38], pc35[38]);
FA1A GS35_39(ps36[38], pc36[39], g35[39], ps35[39], pc35[39]);
FA1A GS35_40(ps36[39], pc36[40], g35[40], ps35[40], pc35[40]);
FA1A GS35_41(ps36[40], pc36[41], g35[41], ps35[41], pc35[41]);
FA1A GS35_42(ps36[41], pc36[42], g35[42], ps35[42], pc35[42]);
FA1A GS35_43(ps36[42], pc36[43], g35[43], ps35[43], pc35[43]);
FA1A GS35_44(ps36[43], pc36[44], g35[44], ps35[44], pc35[44]);
FA1A GS35_45(ps36[44], pc36[45], g35[45], ps35[45], pc35[45]);
FA1A GS35_46(ps36[45], pc36[46], g35[46], ps35[46], pc35[46]);
FA1A GS35_47(ps36[46], pc36[47], g35[47], ps35[47], pc35[47]);
FA1A GS35_48(ps36[47], pc36[48], g35[48], ps35[48], pc35[48]);
FA1A GS35_49(ps36[48], pc36[49], g35[49], ps35[49], pc35[49]);
FA1A GS35_50(ps36[49], pc36[50], g35[50], ps35[50], pc35[50]);
FA1A GS35_51(ps36[50], pc36[51], g35[51], ps35[51], pc35[51]);
FA1A GS35_52(ps36[51], pc36[52], g35[52], ps35[52], pc35[52]);
FA1A GS35_53(ps36[52], pc36[53], g35[53], ps35[53], pc35[53]);
FA1A GS35_54(ps36[53], pc36[54], g35[54], ps35[54], pc35[54]);
FA1A GS35_55(ps36[54], pc36[55], g35[55], ps35[55], pc35[55]);
FA1A GS35_56(ps36[55], pc36[56], g35[56], ps35[56], pc35[56]);
FA1A GS35_57(ps36[56], pc36[57], g35[57], ps35[57], pc35[57]);
FA1A GS35_58(ps36[57], pc36[58], g35[58], ps35[58], pc35[58]);
FA1A GS35_59(ps36[58], pc36[59], g35[59], ps35[59], pc35[59]);
FA1A GS35_60(ps36[59], pc36[60], g35[60], ps35[60], pc35[60]);
FA1A GS35_61(ps36[60], pc36[61], g35[61], ps35[61], pc35[61]);
FA1A GS35_62(ps36[61], pc36[62], g35[62], ps35[62], pc35[62]);
FA1A GS35_63(ps36[62], pc36[63], g35[63], ps35[63], pc35[63]);
FA1A GS34_9(g35[8], pc35[9], g34[9], ps34[9], pc34[9]);
FA1A GS34_10(ps35[9], pc35[10], g34[10], ps34[10], pc34[10]);
FA1A GS34_11(ps35[10], pc35[11], g34[11], ps34[11], pc34[11]);
FA1A GS34_12(ps35[11], pc35[12], g34[12], ps34[12], pc34[12]);
FA1A GS34_13(ps35[12], pc35[13], g34[13], ps34[13], pc34[13]);
FA1A GS34_14(ps35[13], pc35[14], g34[14], ps34[14], pc34[14]);
FA1A GS34_15(ps35[14], pc35[15], g34[15], ps34[15], pc34[15]);
FA1A GS34_16(ps35[15], pc35[16], g34[16], ps34[16], pc34[16]);
FA1A GS34_17(ps35[16], pc35[17], g34[17], ps34[17], pc34[17]);
FA1A GS34_18(ps35[17], pc35[18], g34[18], ps34[18], pc34[18]);
FA1A GS34_19(ps35[18], pc35[19], g34[19], ps34[19], pc34[19]);
FA1A GS34_20(ps35[19], pc35[20], g34[20], ps34[20], pc34[20]);
FA1A GS34_21(ps35[20], pc35[21], g34[21], ps34[21], pc34[21]);
FA1A GS34_22(ps35[21], pc35[22], g34[22], ps34[22], pc34[22]);
FA1A GS34_23(ps35[22], pc35[23], g34[23], ps34[23], pc34[23]);
FA1A GS34_24(ps35[23], pc35[24], g34[24], ps34[24], pc34[24]);
FA1A GS34_25(ps35[24], pc35[25], g34[25], ps34[25], pc34[25]);
FA1A GS34_26(ps35[25], pc35[26], g34[26], ps34[26], pc34[26]);
FA1A GS34_27(ps35[26], pc35[27], g34[27], ps34[27], pc34[27]);
FA1A GS34_28(ps35[27], pc35[28], g34[28], ps34[28], pc34[28]);
FA1A GS34_29(ps35[28], pc35[29], g34[29], ps34[29], pc34[29]);
FA1A GS34_30(ps35[29], pc35[30], g34[30], ps34[30], pc34[30]);
FA1A GS34_31(ps35[30], pc35[31], g34[31], ps34[31], pc34[31]);
FA1A GS34_32(ps35[31], pc35[32], g34[32], ps34[32], pc34[32]);
FA1A GS34_33(ps35[32], pc35[33], g34[33], ps34[33], pc34[33]);
FA1A GS34_34(ps35[33], pc35[34], g34[34], ps34[34], pc34[34]);
FA1A GS34_35(ps35[34], pc35[35], g34[35], ps34[35], pc34[35]);
FA1A GS34_36(ps35[35], pc35[36], g34[36], ps34[36], pc34[36]);
FA1A GS34_37(ps35[36], pc35[37], g34[37], ps34[37], pc34[37]);
FA1A GS34_38(ps35[37], pc35[38], g34[38], ps34[38], pc34[38]);
FA1A GS34_39(ps35[38], pc35[39], g34[39], ps34[39], pc34[39]);
FA1A GS34_40(ps35[39], pc35[40], g34[40], ps34[40], pc34[40]);
FA1A GS34_41(ps35[40], pc35[41], g34[41], ps34[41], pc34[41]);
FA1A GS34_42(ps35[41], pc35[42], g34[42], ps34[42], pc34[42]);
FA1A GS34_43(ps35[42], pc35[43], g34[43], ps34[43], pc34[43]);
FA1A GS34_44(ps35[43], pc35[44], g34[44], ps34[44], pc34[44]);
FA1A GS34_45(ps35[44], pc35[45], g34[45], ps34[45], pc34[45]);
FA1A GS34_46(ps35[45], pc35[46], g34[46], ps34[46], pc34[46]);
FA1A GS34_47(ps35[46], pc35[47], g34[47], ps34[47], pc34[47]);
FA1A GS34_48(ps35[47], pc35[48], g34[48], ps34[48], pc34[48]);
FA1A GS34_49(ps35[48], pc35[49], g34[49], ps34[49], pc34[49]);
FA1A GS34_50(ps35[49], pc35[50], g34[50], ps34[50], pc34[50]);
FA1A GS34_51(ps35[50], pc35[51], g34[51], ps34[51], pc34[51]);
FA1A GS34_52(ps35[51], pc35[52], g34[52], ps34[52], pc34[52]);
FA1A GS34_53(ps35[52], pc35[53], g34[53], ps34[53], pc34[53]);
FA1A GS34_54(ps35[53], pc35[54], g34[54], ps34[54], pc34[54]);
FA1A GS34_55(ps35[54], pc35[55], g34[55], ps34[55], pc34[55]);
FA1A GS34_56(ps35[55], pc35[56], g34[56], ps34[56], pc34[56]);
FA1A GS34_57(ps35[56], pc35[57], g34[57], ps34[57], pc34[57]);
FA1A GS34_58(ps35[57], pc35[58], g34[58], ps34[58], pc34[58]);
FA1A GS34_59(ps35[58], pc35[59], g34[59], ps34[59], pc34[59]);
FA1A GS34_60(ps35[59], pc35[60], g34[60], ps34[60], pc34[60]);
FA1A GS34_61(ps35[60], pc35[61], g34[61], ps34[61], pc34[61]);
FA1A GS34_62(ps35[61], pc35[62], g34[62], ps34[62], pc34[62]);
FA1A GS34_63(ps35[62], pc35[63], g34[63], ps34[63], pc34[63]);
FA1A GS33_9(g34[8], pc34[9], g33[9], ps33[9], pc33[9]);
FA1A GS33_10(ps34[9], pc34[10], g33[10], ps33[10], pc33[10]);
FA1A GS33_11(ps34[10], pc34[11], g33[11], ps33[11], pc33[11]);
FA1A GS33_12(ps34[11], pc34[12], g33[12], ps33[12], pc33[12]);
FA1A GS33_13(ps34[12], pc34[13], g33[13], ps33[13], pc33[13]);
FA1A GS33_14(ps34[13], pc34[14], g33[14], ps33[14], pc33[14]);
FA1A GS33_15(ps34[14], pc34[15], g33[15], ps33[15], pc33[15]);
FA1A GS33_16(ps34[15], pc34[16], g33[16], ps33[16], pc33[16]);
FA1A GS33_17(ps34[16], pc34[17], g33[17], ps33[17], pc33[17]);
FA1A GS33_18(ps34[17], pc34[18], g33[18], ps33[18], pc33[18]);
FA1A GS33_19(ps34[18], pc34[19], g33[19], ps33[19], pc33[19]);
FA1A GS33_20(ps34[19], pc34[20], g33[20], ps33[20], pc33[20]);
FA1A GS33_21(ps34[20], pc34[21], g33[21], ps33[21], pc33[21]);
FA1A GS33_22(ps34[21], pc34[22], g33[22], ps33[22], pc33[22]);
FA1A GS33_23(ps34[22], pc34[23], g33[23], ps33[23], pc33[23]);
FA1A GS33_24(ps34[23], pc34[24], g33[24], ps33[24], pc33[24]);
FA1A GS33_25(ps34[24], pc34[25], g33[25], ps33[25], pc33[25]);
FA1A GS33_26(ps34[25], pc34[26], g33[26], ps33[26], pc33[26]);
FA1A GS33_27(ps34[26], pc34[27], g33[27], ps33[27], pc33[27]);
FA1A GS33_28(ps34[27], pc34[28], g33[28], ps33[28], pc33[28]);
FA1A GS33_29(ps34[28], pc34[29], g33[29], ps33[29], pc33[29]);
FA1A GS33_30(ps34[29], pc34[30], g33[30], ps33[30], pc33[30]);
FA1A GS33_31(ps34[30], pc34[31], g33[31], ps33[31], pc33[31]);
FA1A GS33_32(ps34[31], pc34[32], g33[32], ps33[32], pc33[32]);
FA1A GS33_33(ps34[32], pc34[33], g33[33], ps33[33], pc33[33]);
FA1A GS33_34(ps34[33], pc34[34], g33[34], ps33[34], pc33[34]);
FA1A GS33_35(ps34[34], pc34[35], g33[35], ps33[35], pc33[35]);
FA1A GS33_36(ps34[35], pc34[36], g33[36], ps33[36], pc33[36]);
FA1A GS33_37(ps34[36], pc34[37], g33[37], ps33[37], pc33[37]);
FA1A GS33_38(ps34[37], pc34[38], g33[38], ps33[38], pc33[38]);
FA1A GS33_39(ps34[38], pc34[39], g33[39], ps33[39], pc33[39]);
FA1A GS33_40(ps34[39], pc34[40], g33[40], ps33[40], pc33[40]);
FA1A GS33_41(ps34[40], pc34[41], g33[41], ps33[41], pc33[41]);
FA1A GS33_42(ps34[41], pc34[42], g33[42], ps33[42], pc33[42]);
FA1A GS33_43(ps34[42], pc34[43], g33[43], ps33[43], pc33[43]);
FA1A GS33_44(ps34[43], pc34[44], g33[44], ps33[44], pc33[44]);
FA1A GS33_45(ps34[44], pc34[45], g33[45], ps33[45], pc33[45]);
FA1A GS33_46(ps34[45], pc34[46], g33[46], ps33[46], pc33[46]);
FA1A GS33_47(ps34[46], pc34[47], g33[47], ps33[47], pc33[47]);
FA1A GS33_48(ps34[47], pc34[48], g33[48], ps33[48], pc33[48]);
FA1A GS33_49(ps34[48], pc34[49], g33[49], ps33[49], pc33[49]);
FA1A GS33_50(ps34[49], pc34[50], g33[50], ps33[50], pc33[50]);
FA1A GS33_51(ps34[50], pc34[51], g33[51], ps33[51], pc33[51]);
FA1A GS33_52(ps34[51], pc34[52], g33[52], ps33[52], pc33[52]);
FA1A GS33_53(ps34[52], pc34[53], g33[53], ps33[53], pc33[53]);
FA1A GS33_54(ps34[53], pc34[54], g33[54], ps33[54], pc33[54]);
FA1A GS33_55(ps34[54], pc34[55], g33[55], ps33[55], pc33[55]);
FA1A GS33_56(ps34[55], pc34[56], g33[56], ps33[56], pc33[56]);
FA1A GS33_57(ps34[56], pc34[57], g33[57], ps33[57], pc33[57]);
FA1A GS33_58(ps34[57], pc34[58], g33[58], ps33[58], pc33[58]);
FA1A GS33_59(ps34[58], pc34[59], g33[59], ps33[59], pc33[59]);
FA1A GS33_60(ps34[59], pc34[60], g33[60], ps33[60], pc33[60]);
FA1A GS33_61(ps34[60], pc34[61], g33[61], ps33[61], pc33[61]);
FA1A GS33_62(ps34[61], pc34[62], g33[62], ps33[62], pc33[62]);
FA1A GS33_63(ps34[62], pc34[63], g33[63], ps33[63], pc33[63]);
FA1A GS32_9(g33[8], pc33[9], g32[9], ps32[9], pc32[9]);
FA1A GS32_10(ps33[9], pc33[10], g32[10], ps32[10], pc32[10]);
FA1A GS32_11(ps33[10], pc33[11], g32[11], ps32[11], pc32[11]);
FA1A GS32_12(ps33[11], pc33[12], g32[12], ps32[12], pc32[12]);
FA1A GS32_13(ps33[12], pc33[13], g32[13], ps32[13], pc32[13]);
FA1A GS32_14(ps33[13], pc33[14], g32[14], ps32[14], pc32[14]);
FA1A GS32_15(ps33[14], pc33[15], g32[15], ps32[15], pc32[15]);
FA1A GS32_16(ps33[15], pc33[16], g32[16], ps32[16], pc32[16]);
FA1A GS32_17(ps33[16], pc33[17], g32[17], ps32[17], pc32[17]);
FA1A GS32_18(ps33[17], pc33[18], g32[18], ps32[18], pc32[18]);
FA1A GS32_19(ps33[18], pc33[19], g32[19], ps32[19], pc32[19]);
FA1A GS32_20(ps33[19], pc33[20], g32[20], ps32[20], pc32[20]);
FA1A GS32_21(ps33[20], pc33[21], g32[21], ps32[21], pc32[21]);
FA1A GS32_22(ps33[21], pc33[22], g32[22], ps32[22], pc32[22]);
FA1A GS32_23(ps33[22], pc33[23], g32[23], ps32[23], pc32[23]);
FA1A GS32_24(ps33[23], pc33[24], g32[24], ps32[24], pc32[24]);
FA1A GS32_25(ps33[24], pc33[25], g32[25], ps32[25], pc32[25]);
FA1A GS32_26(ps33[25], pc33[26], g32[26], ps32[26], pc32[26]);
FA1A GS32_27(ps33[26], pc33[27], g32[27], ps32[27], pc32[27]);
FA1A GS32_28(ps33[27], pc33[28], g32[28], ps32[28], pc32[28]);
FA1A GS32_29(ps33[28], pc33[29], g32[29], ps32[29], pc32[29]);
FA1A GS32_30(ps33[29], pc33[30], g32[30], ps32[30], pc32[30]);
FA1A GS32_31(ps33[30], pc33[31], g32[31], ps32[31], pc32[31]);
FA1A GS32_32(ps33[31], pc33[32], g32[32], ps32[32], pc32[32]);
FA1A GS32_33(ps33[32], pc33[33], g32[33], ps32[33], pc32[33]);
FA1A GS32_34(ps33[33], pc33[34], g32[34], ps32[34], pc32[34]);
FA1A GS32_35(ps33[34], pc33[35], g32[35], ps32[35], pc32[35]);
FA1A GS32_36(ps33[35], pc33[36], g32[36], ps32[36], pc32[36]);
FA1A GS32_37(ps33[36], pc33[37], g32[37], ps32[37], pc32[37]);
FA1A GS32_38(ps33[37], pc33[38], g32[38], ps32[38], pc32[38]);
FA1A GS32_39(ps33[38], pc33[39], g32[39], ps32[39], pc32[39]);
FA1A GS32_40(ps33[39], pc33[40], g32[40], ps32[40], pc32[40]);
FA1A GS32_41(ps33[40], pc33[41], g32[41], ps32[41], pc32[41]);
FA1A GS32_42(ps33[41], pc33[42], g32[42], ps32[42], pc32[42]);
FA1A GS32_43(ps33[42], pc33[43], g32[43], ps32[43], pc32[43]);
FA1A GS32_44(ps33[43], pc33[44], g32[44], ps32[44], pc32[44]);
FA1A GS32_45(ps33[44], pc33[45], g32[45], ps32[45], pc32[45]);
FA1A GS32_46(ps33[45], pc33[46], g32[46], ps32[46], pc32[46]);
FA1A GS32_47(ps33[46], pc33[47], g32[47], ps32[47], pc32[47]);
FA1A GS32_48(ps33[47], pc33[48], g32[48], ps32[48], pc32[48]);
FA1A GS32_49(ps33[48], pc33[49], g32[49], ps32[49], pc32[49]);
FA1A GS32_50(ps33[49], pc33[50], g32[50], ps32[50], pc32[50]);
FA1A GS32_51(ps33[50], pc33[51], g32[51], ps32[51], pc32[51]);
FA1A GS32_52(ps33[51], pc33[52], g32[52], ps32[52], pc32[52]);
FA1A GS32_53(ps33[52], pc33[53], g32[53], ps32[53], pc32[53]);
FA1A GS32_54(ps33[53], pc33[54], g32[54], ps32[54], pc32[54]);
FA1A GS32_55(ps33[54], pc33[55], g32[55], ps32[55], pc32[55]);
FA1A GS32_56(ps33[55], pc33[56], g32[56], ps32[56], pc32[56]);
FA1A GS32_57(ps33[56], pc33[57], g32[57], ps32[57], pc32[57]);
FA1A GS32_58(ps33[57], pc33[58], g32[58], ps32[58], pc32[58]);
FA1A GS32_59(ps33[58], pc33[59], g32[59], ps32[59], pc32[59]);
FA1A GS32_60(ps33[59], pc33[60], g32[60], ps32[60], pc32[60]);
FA1A GS32_61(ps33[60], pc33[61], g32[61], ps32[61], pc32[61]);
FA1A GS32_62(ps33[61], pc33[62], g32[62], ps32[62], pc32[62]);
FA1A GS32_63(ps33[62], pc33[63], g32[63], ps32[63], pc32[63]);
FA1A GS31_9(g32[8], pc32[9], g31[9], ps31[9], pc31[9]);
FA1A GS31_10(ps32[9], pc32[10], g31[10], ps31[10], pc31[10]);
FA1A GS31_11(ps32[10], pc32[11], g31[11], ps31[11], pc31[11]);
FA1A GS31_12(ps32[11], pc32[12], g31[12], ps31[12], pc31[12]);
FA1A GS31_13(ps32[12], pc32[13], g31[13], ps31[13], pc31[13]);
FA1A GS31_14(ps32[13], pc32[14], g31[14], ps31[14], pc31[14]);
FA1A GS31_15(ps32[14], pc32[15], g31[15], ps31[15], pc31[15]);
FA1A GS31_16(ps32[15], pc32[16], g31[16], ps31[16], pc31[16]);
FA1A GS31_17(ps32[16], pc32[17], g31[17], ps31[17], pc31[17]);
FA1A GS31_18(ps32[17], pc32[18], g31[18], ps31[18], pc31[18]);
FA1A GS31_19(ps32[18], pc32[19], g31[19], ps31[19], pc31[19]);
FA1A GS31_20(ps32[19], pc32[20], g31[20], ps31[20], pc31[20]);
FA1A GS31_21(ps32[20], pc32[21], g31[21], ps31[21], pc31[21]);
FA1A GS31_22(ps32[21], pc32[22], g31[22], ps31[22], pc31[22]);
FA1A GS31_23(ps32[22], pc32[23], g31[23], ps31[23], pc31[23]);
FA1A GS31_24(ps32[23], pc32[24], g31[24], ps31[24], pc31[24]);
FA1A GS31_25(ps32[24], pc32[25], g31[25], ps31[25], pc31[25]);
FA1A GS31_26(ps32[25], pc32[26], g31[26], ps31[26], pc31[26]);
FA1A GS31_27(ps32[26], pc32[27], g31[27], ps31[27], pc31[27]);
FA1A GS31_28(ps32[27], pc32[28], g31[28], ps31[28], pc31[28]);
FA1A GS31_29(ps32[28], pc32[29], g31[29], ps31[29], pc31[29]);
FA1A GS31_30(ps32[29], pc32[30], g31[30], ps31[30], pc31[30]);
FA1A GS31_31(ps32[30], pc32[31], g31[31], ps31[31], pc31[31]);
FA1A GS31_32(ps32[31], pc32[32], g31[32], ps31[32], pc31[32]);
FA1A GS31_33(ps32[32], pc32[33], g31[33], ps31[33], pc31[33]);
FA1A GS31_34(ps32[33], pc32[34], g31[34], ps31[34], pc31[34]);
FA1A GS31_35(ps32[34], pc32[35], g31[35], ps31[35], pc31[35]);
FA1A GS31_36(ps32[35], pc32[36], g31[36], ps31[36], pc31[36]);
FA1A GS31_37(ps32[36], pc32[37], g31[37], ps31[37], pc31[37]);
FA1A GS31_38(ps32[37], pc32[38], g31[38], ps31[38], pc31[38]);
FA1A GS31_39(ps32[38], pc32[39], g31[39], ps31[39], pc31[39]);
FA1A GS31_40(ps32[39], pc32[40], g31[40], ps31[40], pc31[40]);
FA1A GS31_41(ps32[40], pc32[41], g31[41], ps31[41], pc31[41]);
FA1A GS31_42(ps32[41], pc32[42], g31[42], ps31[42], pc31[42]);
FA1A GS31_43(ps32[42], pc32[43], g31[43], ps31[43], pc31[43]);
FA1A GS31_44(ps32[43], pc32[44], g31[44], ps31[44], pc31[44]);
FA1A GS31_45(ps32[44], pc32[45], g31[45], ps31[45], pc31[45]);
FA1A GS31_46(ps32[45], pc32[46], g31[46], ps31[46], pc31[46]);
FA1A GS31_47(ps32[46], pc32[47], g31[47], ps31[47], pc31[47]);
FA1A GS31_48(ps32[47], pc32[48], g31[48], ps31[48], pc31[48]);
FA1A GS31_49(ps32[48], pc32[49], g31[49], ps31[49], pc31[49]);
FA1A GS31_50(ps32[49], pc32[50], g31[50], ps31[50], pc31[50]);
FA1A GS31_51(ps32[50], pc32[51], g31[51], ps31[51], pc31[51]);
FA1A GS31_52(ps32[51], pc32[52], g31[52], ps31[52], pc31[52]);
FA1A GS31_53(ps32[52], pc32[53], g31[53], ps31[53], pc31[53]);
FA1A GS31_54(ps32[53], pc32[54], g31[54], ps31[54], pc31[54]);
FA1A GS31_55(ps32[54], pc32[55], g31[55], ps31[55], pc31[55]);
FA1A GS31_56(ps32[55], pc32[56], g31[56], ps31[56], pc31[56]);
FA1A GS31_57(ps32[56], pc32[57], g31[57], ps31[57], pc31[57]);
FA1A GS31_58(ps32[57], pc32[58], g31[58], ps31[58], pc31[58]);
FA1A GS31_59(ps32[58], pc32[59], g31[59], ps31[59], pc31[59]);
FA1A GS31_60(ps32[59], pc32[60], g31[60], ps31[60], pc31[60]);
FA1A GS31_61(ps32[60], pc32[61], g31[61], ps31[61], pc31[61]);
FA1A GS31_62(ps32[61], pc32[62], g31[62], ps31[62], pc31[62]);
FA1A GS31_63(ps32[62], pc32[63], g31[63], ps31[63], pc31[63]);
FA1A GS30_9(g31[8], pc31[9], g30[9], ps30[9], pc30[9]);
FA1A GS30_10(ps31[9], pc31[10], g30[10], ps30[10], pc30[10]);
FA1A GS30_11(ps31[10], pc31[11], g30[11], ps30[11], pc30[11]);
FA1A GS30_12(ps31[11], pc31[12], g30[12], ps30[12], pc30[12]);
FA1A GS30_13(ps31[12], pc31[13], g30[13], ps30[13], pc30[13]);
FA1A GS30_14(ps31[13], pc31[14], g30[14], ps30[14], pc30[14]);
FA1A GS30_15(ps31[14], pc31[15], g30[15], ps30[15], pc30[15]);
FA1A GS30_16(ps31[15], pc31[16], g30[16], ps30[16], pc30[16]);
FA1A GS30_17(ps31[16], pc31[17], g30[17], ps30[17], pc30[17]);
FA1A GS30_18(ps31[17], pc31[18], g30[18], ps30[18], pc30[18]);
FA1A GS30_19(ps31[18], pc31[19], g30[19], ps30[19], pc30[19]);
FA1A GS30_20(ps31[19], pc31[20], g30[20], ps30[20], pc30[20]);
FA1A GS30_21(ps31[20], pc31[21], g30[21], ps30[21], pc30[21]);
FA1A GS30_22(ps31[21], pc31[22], g30[22], ps30[22], pc30[22]);
FA1A GS30_23(ps31[22], pc31[23], g30[23], ps30[23], pc30[23]);
FA1A GS30_24(ps31[23], pc31[24], g30[24], ps30[24], pc30[24]);
FA1A GS30_25(ps31[24], pc31[25], g30[25], ps30[25], pc30[25]);
FA1A GS30_26(ps31[25], pc31[26], g30[26], ps30[26], pc30[26]);
FA1A GS30_27(ps31[26], pc31[27], g30[27], ps30[27], pc30[27]);
FA1A GS30_28(ps31[27], pc31[28], g30[28], ps30[28], pc30[28]);
FA1A GS30_29(ps31[28], pc31[29], g30[29], ps30[29], pc30[29]);
FA1A GS30_30(ps31[29], pc31[30], g30[30], ps30[30], pc30[30]);
FA1A GS30_31(ps31[30], pc31[31], g30[31], ps30[31], pc30[31]);
FA1A GS30_32(ps31[31], pc31[32], g30[32], ps30[32], pc30[32]);
FA1A GS30_33(ps31[32], pc31[33], g30[33], ps30[33], pc30[33]);
FA1A GS30_34(ps31[33], pc31[34], g30[34], ps30[34], pc30[34]);
FA1A GS30_35(ps31[34], pc31[35], g30[35], ps30[35], pc30[35]);
FA1A GS30_36(ps31[35], pc31[36], g30[36], ps30[36], pc30[36]);
FA1A GS30_37(ps31[36], pc31[37], g30[37], ps30[37], pc30[37]);
FA1A GS30_38(ps31[37], pc31[38], g30[38], ps30[38], pc30[38]);
FA1A GS30_39(ps31[38], pc31[39], g30[39], ps30[39], pc30[39]);
FA1A GS30_40(ps31[39], pc31[40], g30[40], ps30[40], pc30[40]);
FA1A GS30_41(ps31[40], pc31[41], g30[41], ps30[41], pc30[41]);
FA1A GS30_42(ps31[41], pc31[42], g30[42], ps30[42], pc30[42]);
FA1A GS30_43(ps31[42], pc31[43], g30[43], ps30[43], pc30[43]);
FA1A GS30_44(ps31[43], pc31[44], g30[44], ps30[44], pc30[44]);
FA1A GS30_45(ps31[44], pc31[45], g30[45], ps30[45], pc30[45]);
FA1A GS30_46(ps31[45], pc31[46], g30[46], ps30[46], pc30[46]);
FA1A GS30_47(ps31[46], pc31[47], g30[47], ps30[47], pc30[47]);
FA1A GS30_48(ps31[47], pc31[48], g30[48], ps30[48], pc30[48]);
FA1A GS30_49(ps31[48], pc31[49], g30[49], ps30[49], pc30[49]);
FA1A GS30_50(ps31[49], pc31[50], g30[50], ps30[50], pc30[50]);
FA1A GS30_51(ps31[50], pc31[51], g30[51], ps30[51], pc30[51]);
FA1A GS30_52(ps31[51], pc31[52], g30[52], ps30[52], pc30[52]);
FA1A GS30_53(ps31[52], pc31[53], g30[53], ps30[53], pc30[53]);
FA1A GS30_54(ps31[53], pc31[54], g30[54], ps30[54], pc30[54]);
FA1A GS30_55(ps31[54], pc31[55], g30[55], ps30[55], pc30[55]);
FA1A GS30_56(ps31[55], pc31[56], g30[56], ps30[56], pc30[56]);
FA1A GS30_57(ps31[56], pc31[57], g30[57], ps30[57], pc30[57]);
FA1A GS30_58(ps31[57], pc31[58], g30[58], ps30[58], pc30[58]);
FA1A GS30_59(ps31[58], pc31[59], g30[59], ps30[59], pc30[59]);
FA1A GS30_60(ps31[59], pc31[60], g30[60], ps30[60], pc30[60]);
FA1A GS30_61(ps31[60], pc31[61], g30[61], ps30[61], pc30[61]);
FA1A GS30_62(ps31[61], pc31[62], g30[62], ps30[62], pc30[62]);
FA1A GS30_63(ps31[62], pc31[63], g30[63], ps30[63], pc30[63]);
FA1A GS29_9(g30[8], pc30[9], g29[9], ps29[9], pc29[9]);
FA1A GS29_10(ps30[9], pc30[10], g29[10], ps29[10], pc29[10]);
FA1A GS29_11(ps30[10], pc30[11], g29[11], ps29[11], pc29[11]);
FA1A GS29_12(ps30[11], pc30[12], g29[12], ps29[12], pc29[12]);
FA1A GS29_13(ps30[12], pc30[13], g29[13], ps29[13], pc29[13]);
FA1A GS29_14(ps30[13], pc30[14], g29[14], ps29[14], pc29[14]);
FA1A GS29_15(ps30[14], pc30[15], g29[15], ps29[15], pc29[15]);
FA1A GS29_16(ps30[15], pc30[16], g29[16], ps29[16], pc29[16]);
FA1A GS29_17(ps30[16], pc30[17], g29[17], ps29[17], pc29[17]);
FA1A GS29_18(ps30[17], pc30[18], g29[18], ps29[18], pc29[18]);
FA1A GS29_19(ps30[18], pc30[19], g29[19], ps29[19], pc29[19]);
FA1A GS29_20(ps30[19], pc30[20], g29[20], ps29[20], pc29[20]);
FA1A GS29_21(ps30[20], pc30[21], g29[21], ps29[21], pc29[21]);
FA1A GS29_22(ps30[21], pc30[22], g29[22], ps29[22], pc29[22]);
FA1A GS29_23(ps30[22], pc30[23], g29[23], ps29[23], pc29[23]);
FA1A GS29_24(ps30[23], pc30[24], g29[24], ps29[24], pc29[24]);
FA1A GS29_25(ps30[24], pc30[25], g29[25], ps29[25], pc29[25]);
FA1A GS29_26(ps30[25], pc30[26], g29[26], ps29[26], pc29[26]);
FA1A GS29_27(ps30[26], pc30[27], g29[27], ps29[27], pc29[27]);
FA1A GS29_28(ps30[27], pc30[28], g29[28], ps29[28], pc29[28]);
FA1A GS29_29(ps30[28], pc30[29], g29[29], ps29[29], pc29[29]);
FA1A GS29_30(ps30[29], pc30[30], g29[30], ps29[30], pc29[30]);
FA1A GS29_31(ps30[30], pc30[31], g29[31], ps29[31], pc29[31]);
FA1A GS29_32(ps30[31], pc30[32], g29[32], ps29[32], pc29[32]);
FA1A GS29_33(ps30[32], pc30[33], g29[33], ps29[33], pc29[33]);
FA1A GS29_34(ps30[33], pc30[34], g29[34], ps29[34], pc29[34]);
FA1A GS29_35(ps30[34], pc30[35], g29[35], ps29[35], pc29[35]);
FA1A GS29_36(ps30[35], pc30[36], g29[36], ps29[36], pc29[36]);
FA1A GS29_37(ps30[36], pc30[37], g29[37], ps29[37], pc29[37]);
FA1A GS29_38(ps30[37], pc30[38], g29[38], ps29[38], pc29[38]);
FA1A GS29_39(ps30[38], pc30[39], g29[39], ps29[39], pc29[39]);
FA1A GS29_40(ps30[39], pc30[40], g29[40], ps29[40], pc29[40]);
FA1A GS29_41(ps30[40], pc30[41], g29[41], ps29[41], pc29[41]);
FA1A GS29_42(ps30[41], pc30[42], g29[42], ps29[42], pc29[42]);
FA1A GS29_43(ps30[42], pc30[43], g29[43], ps29[43], pc29[43]);
FA1A GS29_44(ps30[43], pc30[44], g29[44], ps29[44], pc29[44]);
FA1A GS29_45(ps30[44], pc30[45], g29[45], ps29[45], pc29[45]);
FA1A GS29_46(ps30[45], pc30[46], g29[46], ps29[46], pc29[46]);
FA1A GS29_47(ps30[46], pc30[47], g29[47], ps29[47], pc29[47]);
FA1A GS29_48(ps30[47], pc30[48], g29[48], ps29[48], pc29[48]);
FA1A GS29_49(ps30[48], pc30[49], g29[49], ps29[49], pc29[49]);
FA1A GS29_50(ps30[49], pc30[50], g29[50], ps29[50], pc29[50]);
FA1A GS29_51(ps30[50], pc30[51], g29[51], ps29[51], pc29[51]);
FA1A GS29_52(ps30[51], pc30[52], g29[52], ps29[52], pc29[52]);
FA1A GS29_53(ps30[52], pc30[53], g29[53], ps29[53], pc29[53]);
FA1A GS29_54(ps30[53], pc30[54], g29[54], ps29[54], pc29[54]);
FA1A GS29_55(ps30[54], pc30[55], g29[55], ps29[55], pc29[55]);
FA1A GS29_56(ps30[55], pc30[56], g29[56], ps29[56], pc29[56]);
FA1A GS29_57(ps30[56], pc30[57], g29[57], ps29[57], pc29[57]);
FA1A GS29_58(ps30[57], pc30[58], g29[58], ps29[58], pc29[58]);
FA1A GS29_59(ps30[58], pc30[59], g29[59], ps29[59], pc29[59]);
FA1A GS29_60(ps30[59], pc30[60], g29[60], ps29[60], pc29[60]);
FA1A GS29_61(ps30[60], pc30[61], g29[61], ps29[61], pc29[61]);
FA1A GS29_62(ps30[61], pc30[62], g29[62], ps29[62], pc29[62]);
FA1A GS29_63(ps30[62], pc30[63], g29[63], ps29[63], pc29[63]);
FA1A GS28_9(g29[8], pc29[9], g28[9], ps28[9], pc28[9]);
FA1A GS28_10(ps29[9], pc29[10], g28[10], ps28[10], pc28[10]);
FA1A GS28_11(ps29[10], pc29[11], g28[11], ps28[11], pc28[11]);
FA1A GS28_12(ps29[11], pc29[12], g28[12], ps28[12], pc28[12]);
FA1A GS28_13(ps29[12], pc29[13], g28[13], ps28[13], pc28[13]);
FA1A GS28_14(ps29[13], pc29[14], g28[14], ps28[14], pc28[14]);
FA1A GS28_15(ps29[14], pc29[15], g28[15], ps28[15], pc28[15]);
FA1A GS28_16(ps29[15], pc29[16], g28[16], ps28[16], pc28[16]);
FA1A GS28_17(ps29[16], pc29[17], g28[17], ps28[17], pc28[17]);
FA1A GS28_18(ps29[17], pc29[18], g28[18], ps28[18], pc28[18]);
FA1A GS28_19(ps29[18], pc29[19], g28[19], ps28[19], pc28[19]);
FA1A GS28_20(ps29[19], pc29[20], g28[20], ps28[20], pc28[20]);
FA1A GS28_21(ps29[20], pc29[21], g28[21], ps28[21], pc28[21]);
FA1A GS28_22(ps29[21], pc29[22], g28[22], ps28[22], pc28[22]);
FA1A GS28_23(ps29[22], pc29[23], g28[23], ps28[23], pc28[23]);
FA1A GS28_24(ps29[23], pc29[24], g28[24], ps28[24], pc28[24]);
FA1A GS28_25(ps29[24], pc29[25], g28[25], ps28[25], pc28[25]);
FA1A GS28_26(ps29[25], pc29[26], g28[26], ps28[26], pc28[26]);
FA1A GS28_27(ps29[26], pc29[27], g28[27], ps28[27], pc28[27]);
FA1A GS28_28(ps29[27], pc29[28], g28[28], ps28[28], pc28[28]);
FA1A GS28_29(ps29[28], pc29[29], g28[29], ps28[29], pc28[29]);
FA1A GS28_30(ps29[29], pc29[30], g28[30], ps28[30], pc28[30]);
FA1A GS28_31(ps29[30], pc29[31], g28[31], ps28[31], pc28[31]);
FA1A GS28_32(ps29[31], pc29[32], g28[32], ps28[32], pc28[32]);
FA1A GS28_33(ps29[32], pc29[33], g28[33], ps28[33], pc28[33]);
FA1A GS28_34(ps29[33], pc29[34], g28[34], ps28[34], pc28[34]);
FA1A GS28_35(ps29[34], pc29[35], g28[35], ps28[35], pc28[35]);
FA1A GS28_36(ps29[35], pc29[36], g28[36], ps28[36], pc28[36]);
FA1A GS28_37(ps29[36], pc29[37], g28[37], ps28[37], pc28[37]);
FA1A GS28_38(ps29[37], pc29[38], g28[38], ps28[38], pc28[38]);
FA1A GS28_39(ps29[38], pc29[39], g28[39], ps28[39], pc28[39]);
FA1A GS28_40(ps29[39], pc29[40], g28[40], ps28[40], pc28[40]);
FA1A GS28_41(ps29[40], pc29[41], g28[41], ps28[41], pc28[41]);
FA1A GS28_42(ps29[41], pc29[42], g28[42], ps28[42], pc28[42]);
FA1A GS28_43(ps29[42], pc29[43], g28[43], ps28[43], pc28[43]);
FA1A GS28_44(ps29[43], pc29[44], g28[44], ps28[44], pc28[44]);
FA1A GS28_45(ps29[44], pc29[45], g28[45], ps28[45], pc28[45]);
FA1A GS28_46(ps29[45], pc29[46], g28[46], ps28[46], pc28[46]);
FA1A GS28_47(ps29[46], pc29[47], g28[47], ps28[47], pc28[47]);
FA1A GS28_48(ps29[47], pc29[48], g28[48], ps28[48], pc28[48]);
FA1A GS28_49(ps29[48], pc29[49], g28[49], ps28[49], pc28[49]);
FA1A GS28_50(ps29[49], pc29[50], g28[50], ps28[50], pc28[50]);
FA1A GS28_51(ps29[50], pc29[51], g28[51], ps28[51], pc28[51]);
FA1A GS28_52(ps29[51], pc29[52], g28[52], ps28[52], pc28[52]);
FA1A GS28_53(ps29[52], pc29[53], g28[53], ps28[53], pc28[53]);
FA1A GS28_54(ps29[53], pc29[54], g28[54], ps28[54], pc28[54]);
FA1A GS28_55(ps29[54], pc29[55], g28[55], ps28[55], pc28[55]);
FA1A GS28_56(ps29[55], pc29[56], g28[56], ps28[56], pc28[56]);
FA1A GS28_57(ps29[56], pc29[57], g28[57], ps28[57], pc28[57]);
FA1A GS28_58(ps29[57], pc29[58], g28[58], ps28[58], pc28[58]);
FA1A GS28_59(ps29[58], pc29[59], g28[59], ps28[59], pc28[59]);
FA1A GS28_60(ps29[59], pc29[60], g28[60], ps28[60], pc28[60]);
FA1A GS28_61(ps29[60], pc29[61], g28[61], ps28[61], pc28[61]);
FA1A GS28_62(ps29[61], pc29[62], g28[62], ps28[62], pc28[62]);
FA1A GS28_63(ps29[62], pc29[63], g28[63], ps28[63], pc28[63]);
FA1A GS27_9(g28[8], pc28[9], g27[9], ps27[9], pc27[9]);
FA1A GS27_10(ps28[9], pc28[10], g27[10], ps27[10], pc27[10]);
FA1A GS27_11(ps28[10], pc28[11], g27[11], ps27[11], pc27[11]);
FA1A GS27_12(ps28[11], pc28[12], g27[12], ps27[12], pc27[12]);
FA1A GS27_13(ps28[12], pc28[13], g27[13], ps27[13], pc27[13]);
FA1A GS27_14(ps28[13], pc28[14], g27[14], ps27[14], pc27[14]);
FA1A GS27_15(ps28[14], pc28[15], g27[15], ps27[15], pc27[15]);
FA1A GS27_16(ps28[15], pc28[16], g27[16], ps27[16], pc27[16]);
FA1A GS27_17(ps28[16], pc28[17], g27[17], ps27[17], pc27[17]);
FA1A GS27_18(ps28[17], pc28[18], g27[18], ps27[18], pc27[18]);
FA1A GS27_19(ps28[18], pc28[19], g27[19], ps27[19], pc27[19]);
FA1A GS27_20(ps28[19], pc28[20], g27[20], ps27[20], pc27[20]);
FA1A GS27_21(ps28[20], pc28[21], g27[21], ps27[21], pc27[21]);
FA1A GS27_22(ps28[21], pc28[22], g27[22], ps27[22], pc27[22]);
FA1A GS27_23(ps28[22], pc28[23], g27[23], ps27[23], pc27[23]);
FA1A GS27_24(ps28[23], pc28[24], g27[24], ps27[24], pc27[24]);
FA1A GS27_25(ps28[24], pc28[25], g27[25], ps27[25], pc27[25]);
FA1A GS27_26(ps28[25], pc28[26], g27[26], ps27[26], pc27[26]);
FA1A GS27_27(ps28[26], pc28[27], g27[27], ps27[27], pc27[27]);
FA1A GS27_28(ps28[27], pc28[28], g27[28], ps27[28], pc27[28]);
FA1A GS27_29(ps28[28], pc28[29], g27[29], ps27[29], pc27[29]);
FA1A GS27_30(ps28[29], pc28[30], g27[30], ps27[30], pc27[30]);
FA1A GS27_31(ps28[30], pc28[31], g27[31], ps27[31], pc27[31]);
FA1A GS27_32(ps28[31], pc28[32], g27[32], ps27[32], pc27[32]);
FA1A GS27_33(ps28[32], pc28[33], g27[33], ps27[33], pc27[33]);
FA1A GS27_34(ps28[33], pc28[34], g27[34], ps27[34], pc27[34]);
FA1A GS27_35(ps28[34], pc28[35], g27[35], ps27[35], pc27[35]);
FA1A GS27_36(ps28[35], pc28[36], g27[36], ps27[36], pc27[36]);
FA1A GS27_37(ps28[36], pc28[37], g27[37], ps27[37], pc27[37]);
FA1A GS27_38(ps28[37], pc28[38], g27[38], ps27[38], pc27[38]);
FA1A GS27_39(ps28[38], pc28[39], g27[39], ps27[39], pc27[39]);
FA1A GS27_40(ps28[39], pc28[40], g27[40], ps27[40], pc27[40]);
FA1A GS27_41(ps28[40], pc28[41], g27[41], ps27[41], pc27[41]);
FA1A GS27_42(ps28[41], pc28[42], g27[42], ps27[42], pc27[42]);
FA1A GS27_43(ps28[42], pc28[43], g27[43], ps27[43], pc27[43]);
FA1A GS27_44(ps28[43], pc28[44], g27[44], ps27[44], pc27[44]);
FA1A GS27_45(ps28[44], pc28[45], g27[45], ps27[45], pc27[45]);
FA1A GS27_46(ps28[45], pc28[46], g27[46], ps27[46], pc27[46]);
FA1A GS27_47(ps28[46], pc28[47], g27[47], ps27[47], pc27[47]);
FA1A GS27_48(ps28[47], pc28[48], g27[48], ps27[48], pc27[48]);
FA1A GS27_49(ps28[48], pc28[49], g27[49], ps27[49], pc27[49]);
FA1A GS27_50(ps28[49], pc28[50], g27[50], ps27[50], pc27[50]);
FA1A GS27_51(ps28[50], pc28[51], g27[51], ps27[51], pc27[51]);
FA1A GS27_52(ps28[51], pc28[52], g27[52], ps27[52], pc27[52]);
FA1A GS27_53(ps28[52], pc28[53], g27[53], ps27[53], pc27[53]);
FA1A GS27_54(ps28[53], pc28[54], g27[54], ps27[54], pc27[54]);
FA1A GS27_55(ps28[54], pc28[55], g27[55], ps27[55], pc27[55]);
FA1A GS27_56(ps28[55], pc28[56], g27[56], ps27[56], pc27[56]);
FA1A GS27_57(ps28[56], pc28[57], g27[57], ps27[57], pc27[57]);
FA1A GS27_58(ps28[57], pc28[58], g27[58], ps27[58], pc27[58]);
FA1A GS27_59(ps28[58], pc28[59], g27[59], ps27[59], pc27[59]);
FA1A GS27_60(ps28[59], pc28[60], g27[60], ps27[60], pc27[60]);
FA1A GS27_61(ps28[60], pc28[61], g27[61], ps27[61], pc27[61]);
FA1A GS27_62(ps28[61], pc28[62], g27[62], ps27[62], pc27[62]);
FA1A GS27_63(ps28[62], pc28[63], g27[63], ps27[63], pc27[63]);
FA1A GS26_9(g27[8], pc27[9], g26[9], ps26[9], pc26[9]);
FA1A GS26_10(ps27[9], pc27[10], g26[10], ps26[10], pc26[10]);
FA1A GS26_11(ps27[10], pc27[11], g26[11], ps26[11], pc26[11]);
FA1A GS26_12(ps27[11], pc27[12], g26[12], ps26[12], pc26[12]);
FA1A GS26_13(ps27[12], pc27[13], g26[13], ps26[13], pc26[13]);
FA1A GS26_14(ps27[13], pc27[14], g26[14], ps26[14], pc26[14]);
FA1A GS26_15(ps27[14], pc27[15], g26[15], ps26[15], pc26[15]);
FA1A GS26_16(ps27[15], pc27[16], g26[16], ps26[16], pc26[16]);
FA1A GS26_17(ps27[16], pc27[17], g26[17], ps26[17], pc26[17]);
FA1A GS26_18(ps27[17], pc27[18], g26[18], ps26[18], pc26[18]);
FA1A GS26_19(ps27[18], pc27[19], g26[19], ps26[19], pc26[19]);
FA1A GS26_20(ps27[19], pc27[20], g26[20], ps26[20], pc26[20]);
FA1A GS26_21(ps27[20], pc27[21], g26[21], ps26[21], pc26[21]);
FA1A GS26_22(ps27[21], pc27[22], g26[22], ps26[22], pc26[22]);
FA1A GS26_23(ps27[22], pc27[23], g26[23], ps26[23], pc26[23]);
FA1A GS26_24(ps27[23], pc27[24], g26[24], ps26[24], pc26[24]);
FA1A GS26_25(ps27[24], pc27[25], g26[25], ps26[25], pc26[25]);
FA1A GS26_26(ps27[25], pc27[26], g26[26], ps26[26], pc26[26]);
FA1A GS26_27(ps27[26], pc27[27], g26[27], ps26[27], pc26[27]);
FA1A GS26_28(ps27[27], pc27[28], g26[28], ps26[28], pc26[28]);
FA1A GS26_29(ps27[28], pc27[29], g26[29], ps26[29], pc26[29]);
FA1A GS26_30(ps27[29], pc27[30], g26[30], ps26[30], pc26[30]);
FA1A GS26_31(ps27[30], pc27[31], g26[31], ps26[31], pc26[31]);
FA1A GS26_32(ps27[31], pc27[32], g26[32], ps26[32], pc26[32]);
FA1A GS26_33(ps27[32], pc27[33], g26[33], ps26[33], pc26[33]);
FA1A GS26_34(ps27[33], pc27[34], g26[34], ps26[34], pc26[34]);
FA1A GS26_35(ps27[34], pc27[35], g26[35], ps26[35], pc26[35]);
FA1A GS26_36(ps27[35], pc27[36], g26[36], ps26[36], pc26[36]);
FA1A GS26_37(ps27[36], pc27[37], g26[37], ps26[37], pc26[37]);
FA1A GS26_38(ps27[37], pc27[38], g26[38], ps26[38], pc26[38]);
FA1A GS26_39(ps27[38], pc27[39], g26[39], ps26[39], pc26[39]);
FA1A GS26_40(ps27[39], pc27[40], g26[40], ps26[40], pc26[40]);
FA1A GS26_41(ps27[40], pc27[41], g26[41], ps26[41], pc26[41]);
FA1A GS26_42(ps27[41], pc27[42], g26[42], ps26[42], pc26[42]);
FA1A GS26_43(ps27[42], pc27[43], g26[43], ps26[43], pc26[43]);
FA1A GS26_44(ps27[43], pc27[44], g26[44], ps26[44], pc26[44]);
FA1A GS26_45(ps27[44], pc27[45], g26[45], ps26[45], pc26[45]);
FA1A GS26_46(ps27[45], pc27[46], g26[46], ps26[46], pc26[46]);
FA1A GS26_47(ps27[46], pc27[47], g26[47], ps26[47], pc26[47]);
FA1A GS26_48(ps27[47], pc27[48], g26[48], ps26[48], pc26[48]);
FA1A GS26_49(ps27[48], pc27[49], g26[49], ps26[49], pc26[49]);
FA1A GS26_50(ps27[49], pc27[50], g26[50], ps26[50], pc26[50]);
FA1A GS26_51(ps27[50], pc27[51], g26[51], ps26[51], pc26[51]);
FA1A GS26_52(ps27[51], pc27[52], g26[52], ps26[52], pc26[52]);
FA1A GS26_53(ps27[52], pc27[53], g26[53], ps26[53], pc26[53]);
FA1A GS26_54(ps27[53], pc27[54], g26[54], ps26[54], pc26[54]);
FA1A GS26_55(ps27[54], pc27[55], g26[55], ps26[55], pc26[55]);
FA1A GS26_56(ps27[55], pc27[56], g26[56], ps26[56], pc26[56]);
FA1A GS26_57(ps27[56], pc27[57], g26[57], ps26[57], pc26[57]);
FA1A GS26_58(ps27[57], pc27[58], g26[58], ps26[58], pc26[58]);
FA1A GS26_59(ps27[58], pc27[59], g26[59], ps26[59], pc26[59]);
FA1A GS26_60(ps27[59], pc27[60], g26[60], ps26[60], pc26[60]);
FA1A GS26_61(ps27[60], pc27[61], g26[61], ps26[61], pc26[61]);
FA1A GS26_62(ps27[61], pc27[62], g26[62], ps26[62], pc26[62]);
FA1A GS26_63(ps27[62], pc27[63], g26[63], ps26[63], pc26[63]);
FA1A GS25_9(g26[8], pc26[9], g25[9], ps25[9], pc25[9]);
FA1A GS25_10(ps26[9], pc26[10], g25[10], ps25[10], pc25[10]);
FA1A GS25_11(ps26[10], pc26[11], g25[11], ps25[11], pc25[11]);
FA1A GS25_12(ps26[11], pc26[12], g25[12], ps25[12], pc25[12]);
FA1A GS25_13(ps26[12], pc26[13], g25[13], ps25[13], pc25[13]);
FA1A GS25_14(ps26[13], pc26[14], g25[14], ps25[14], pc25[14]);
FA1A GS25_15(ps26[14], pc26[15], g25[15], ps25[15], pc25[15]);
FA1A GS25_16(ps26[15], pc26[16], g25[16], ps25[16], pc25[16]);
FA1A GS25_17(ps26[16], pc26[17], g25[17], ps25[17], pc25[17]);
FA1A GS25_18(ps26[17], pc26[18], g25[18], ps25[18], pc25[18]);
FA1A GS25_19(ps26[18], pc26[19], g25[19], ps25[19], pc25[19]);
FA1A GS25_20(ps26[19], pc26[20], g25[20], ps25[20], pc25[20]);
FA1A GS25_21(ps26[20], pc26[21], g25[21], ps25[21], pc25[21]);
FA1A GS25_22(ps26[21], pc26[22], g25[22], ps25[22], pc25[22]);
FA1A GS25_23(ps26[22], pc26[23], g25[23], ps25[23], pc25[23]);
FA1A GS25_24(ps26[23], pc26[24], g25[24], ps25[24], pc25[24]);
FA1A GS25_25(ps26[24], pc26[25], g25[25], ps25[25], pc25[25]);
FA1A GS25_26(ps26[25], pc26[26], g25[26], ps25[26], pc25[26]);
FA1A GS25_27(ps26[26], pc26[27], g25[27], ps25[27], pc25[27]);
FA1A GS25_28(ps26[27], pc26[28], g25[28], ps25[28], pc25[28]);
FA1A GS25_29(ps26[28], pc26[29], g25[29], ps25[29], pc25[29]);
FA1A GS25_30(ps26[29], pc26[30], g25[30], ps25[30], pc25[30]);
FA1A GS25_31(ps26[30], pc26[31], g25[31], ps25[31], pc25[31]);
FA1A GS25_32(ps26[31], pc26[32], g25[32], ps25[32], pc25[32]);
FA1A GS25_33(ps26[32], pc26[33], g25[33], ps25[33], pc25[33]);
FA1A GS25_34(ps26[33], pc26[34], g25[34], ps25[34], pc25[34]);
FA1A GS25_35(ps26[34], pc26[35], g25[35], ps25[35], pc25[35]);
FA1A GS25_36(ps26[35], pc26[36], g25[36], ps25[36], pc25[36]);
FA1A GS25_37(ps26[36], pc26[37], g25[37], ps25[37], pc25[37]);
FA1A GS25_38(ps26[37], pc26[38], g25[38], ps25[38], pc25[38]);
FA1A GS25_39(ps26[38], pc26[39], g25[39], ps25[39], pc25[39]);
FA1A GS25_40(ps26[39], pc26[40], g25[40], ps25[40], pc25[40]);
FA1A GS25_41(ps26[40], pc26[41], g25[41], ps25[41], pc25[41]);
FA1A GS25_42(ps26[41], pc26[42], g25[42], ps25[42], pc25[42]);
FA1A GS25_43(ps26[42], pc26[43], g25[43], ps25[43], pc25[43]);
FA1A GS25_44(ps26[43], pc26[44], g25[44], ps25[44], pc25[44]);
FA1A GS25_45(ps26[44], pc26[45], g25[45], ps25[45], pc25[45]);
FA1A GS25_46(ps26[45], pc26[46], g25[46], ps25[46], pc25[46]);
FA1A GS25_47(ps26[46], pc26[47], g25[47], ps25[47], pc25[47]);
FA1A GS25_48(ps26[47], pc26[48], g25[48], ps25[48], pc25[48]);
FA1A GS25_49(ps26[48], pc26[49], g25[49], ps25[49], pc25[49]);
FA1A GS25_50(ps26[49], pc26[50], g25[50], ps25[50], pc25[50]);
FA1A GS25_51(ps26[50], pc26[51], g25[51], ps25[51], pc25[51]);
FA1A GS25_52(ps26[51], pc26[52], g25[52], ps25[52], pc25[52]);
FA1A GS25_53(ps26[52], pc26[53], g25[53], ps25[53], pc25[53]);
FA1A GS25_54(ps26[53], pc26[54], g25[54], ps25[54], pc25[54]);
FA1A GS25_55(ps26[54], pc26[55], g25[55], ps25[55], pc25[55]);
FA1A GS25_56(ps26[55], pc26[56], g25[56], ps25[56], pc25[56]);
FA1A GS25_57(ps26[56], pc26[57], g25[57], ps25[57], pc25[57]);
FA1A GS25_58(ps26[57], pc26[58], g25[58], ps25[58], pc25[58]);
FA1A GS25_59(ps26[58], pc26[59], g25[59], ps25[59], pc25[59]);
FA1A GS25_60(ps26[59], pc26[60], g25[60], ps25[60], pc25[60]);
FA1A GS25_61(ps26[60], pc26[61], g25[61], ps25[61], pc25[61]);
FA1A GS25_62(ps26[61], pc26[62], g25[62], ps25[62], pc25[62]);
FA1A GS25_63(ps26[62], pc26[63], g25[63], ps25[63], pc25[63]);
FA1A GS24_9(g25[8], pc25[9], g24[9], ps24[9], pc24[9]);
FA1A GS24_10(ps25[9], pc25[10], g24[10], ps24[10], pc24[10]);
FA1A GS24_11(ps25[10], pc25[11], g24[11], ps24[11], pc24[11]);
FA1A GS24_12(ps25[11], pc25[12], g24[12], ps24[12], pc24[12]);
FA1A GS24_13(ps25[12], pc25[13], g24[13], ps24[13], pc24[13]);
FA1A GS24_14(ps25[13], pc25[14], g24[14], ps24[14], pc24[14]);
FA1A GS24_15(ps25[14], pc25[15], g24[15], ps24[15], pc24[15]);
FA1A GS24_16(ps25[15], pc25[16], g24[16], ps24[16], pc24[16]);
FA1A GS24_17(ps25[16], pc25[17], g24[17], ps24[17], pc24[17]);
FA1A GS24_18(ps25[17], pc25[18], g24[18], ps24[18], pc24[18]);
FA1A GS24_19(ps25[18], pc25[19], g24[19], ps24[19], pc24[19]);
FA1A GS24_20(ps25[19], pc25[20], g24[20], ps24[20], pc24[20]);
FA1A GS24_21(ps25[20], pc25[21], g24[21], ps24[21], pc24[21]);
FA1A GS24_22(ps25[21], pc25[22], g24[22], ps24[22], pc24[22]);
FA1A GS24_23(ps25[22], pc25[23], g24[23], ps24[23], pc24[23]);
FA1A GS24_24(ps25[23], pc25[24], g24[24], ps24[24], pc24[24]);
FA1A GS24_25(ps25[24], pc25[25], g24[25], ps24[25], pc24[25]);
FA1A GS24_26(ps25[25], pc25[26], g24[26], ps24[26], pc24[26]);
FA1A GS24_27(ps25[26], pc25[27], g24[27], ps24[27], pc24[27]);
FA1A GS24_28(ps25[27], pc25[28], g24[28], ps24[28], pc24[28]);
FA1A GS24_29(ps25[28], pc25[29], g24[29], ps24[29], pc24[29]);
FA1A GS24_30(ps25[29], pc25[30], g24[30], ps24[30], pc24[30]);
FA1A GS24_31(ps25[30], pc25[31], g24[31], ps24[31], pc24[31]);
FA1A GS24_32(ps25[31], pc25[32], g24[32], ps24[32], pc24[32]);
FA1A GS24_33(ps25[32], pc25[33], g24[33], ps24[33], pc24[33]);
FA1A GS24_34(ps25[33], pc25[34], g24[34], ps24[34], pc24[34]);
FA1A GS24_35(ps25[34], pc25[35], g24[35], ps24[35], pc24[35]);
FA1A GS24_36(ps25[35], pc25[36], g24[36], ps24[36], pc24[36]);
FA1A GS24_37(ps25[36], pc25[37], g24[37], ps24[37], pc24[37]);
FA1A GS24_38(ps25[37], pc25[38], g24[38], ps24[38], pc24[38]);
FA1A GS24_39(ps25[38], pc25[39], g24[39], ps24[39], pc24[39]);
FA1A GS24_40(ps25[39], pc25[40], g24[40], ps24[40], pc24[40]);
FA1A GS24_41(ps25[40], pc25[41], g24[41], ps24[41], pc24[41]);
FA1A GS24_42(ps25[41], pc25[42], g24[42], ps24[42], pc24[42]);
FA1A GS24_43(ps25[42], pc25[43], g24[43], ps24[43], pc24[43]);
FA1A GS24_44(ps25[43], pc25[44], g24[44], ps24[44], pc24[44]);
FA1A GS24_45(ps25[44], pc25[45], g24[45], ps24[45], pc24[45]);
FA1A GS24_46(ps25[45], pc25[46], g24[46], ps24[46], pc24[46]);
FA1A GS24_47(ps25[46], pc25[47], g24[47], ps24[47], pc24[47]);
FA1A GS24_48(ps25[47], pc25[48], g24[48], ps24[48], pc24[48]);
FA1A GS24_49(ps25[48], pc25[49], g24[49], ps24[49], pc24[49]);
FA1A GS24_50(ps25[49], pc25[50], g24[50], ps24[50], pc24[50]);
FA1A GS24_51(ps25[50], pc25[51], g24[51], ps24[51], pc24[51]);
FA1A GS24_52(ps25[51], pc25[52], g24[52], ps24[52], pc24[52]);
FA1A GS24_53(ps25[52], pc25[53], g24[53], ps24[53], pc24[53]);
FA1A GS24_54(ps25[53], pc25[54], g24[54], ps24[54], pc24[54]);
FA1A GS24_55(ps25[54], pc25[55], g24[55], ps24[55], pc24[55]);
FA1A GS24_56(ps25[55], pc25[56], g24[56], ps24[56], pc24[56]);
FA1A GS24_57(ps25[56], pc25[57], g24[57], ps24[57], pc24[57]);
FA1A GS24_58(ps25[57], pc25[58], g24[58], ps24[58], pc24[58]);
FA1A GS24_59(ps25[58], pc25[59], g24[59], ps24[59], pc24[59]);
FA1A GS24_60(ps25[59], pc25[60], g24[60], ps24[60], pc24[60]);
FA1A GS24_61(ps25[60], pc25[61], g24[61], ps24[61], pc24[61]);
FA1A GS24_62(ps25[61], pc25[62], g24[62], ps24[62], pc24[62]);
FA1A GS24_63(ps25[62], pc25[63], g24[63], ps24[63], pc24[63]);
FA1A GS23_9(g24[8], pc24[9], g23[9], ps23[9], pc23[9]);
FA1A GS23_10(ps24[9], pc24[10], g23[10], ps23[10], pc23[10]);
FA1A GS23_11(ps24[10], pc24[11], g23[11], ps23[11], pc23[11]);
FA1A GS23_12(ps24[11], pc24[12], g23[12], ps23[12], pc23[12]);
FA1A GS23_13(ps24[12], pc24[13], g23[13], ps23[13], pc23[13]);
FA1A GS23_14(ps24[13], pc24[14], g23[14], ps23[14], pc23[14]);
FA1A GS23_15(ps24[14], pc24[15], g23[15], ps23[15], pc23[15]);
FA1A GS23_16(ps24[15], pc24[16], g23[16], ps23[16], pc23[16]);
FA1A GS23_17(ps24[16], pc24[17], g23[17], ps23[17], pc23[17]);
FA1A GS23_18(ps24[17], pc24[18], g23[18], ps23[18], pc23[18]);
FA1A GS23_19(ps24[18], pc24[19], g23[19], ps23[19], pc23[19]);
FA1A GS23_20(ps24[19], pc24[20], g23[20], ps23[20], pc23[20]);
FA1A GS23_21(ps24[20], pc24[21], g23[21], ps23[21], pc23[21]);
FA1A GS23_22(ps24[21], pc24[22], g23[22], ps23[22], pc23[22]);
FA1A GS23_23(ps24[22], pc24[23], g23[23], ps23[23], pc23[23]);
FA1A GS23_24(ps24[23], pc24[24], g23[24], ps23[24], pc23[24]);
FA1A GS23_25(ps24[24], pc24[25], g23[25], ps23[25], pc23[25]);
FA1A GS23_26(ps24[25], pc24[26], g23[26], ps23[26], pc23[26]);
FA1A GS23_27(ps24[26], pc24[27], g23[27], ps23[27], pc23[27]);
FA1A GS23_28(ps24[27], pc24[28], g23[28], ps23[28], pc23[28]);
FA1A GS23_29(ps24[28], pc24[29], g23[29], ps23[29], pc23[29]);
FA1A GS23_30(ps24[29], pc24[30], g23[30], ps23[30], pc23[30]);
FA1A GS23_31(ps24[30], pc24[31], g23[31], ps23[31], pc23[31]);
FA1A GS23_32(ps24[31], pc24[32], g23[32], ps23[32], pc23[32]);
FA1A GS23_33(ps24[32], pc24[33], g23[33], ps23[33], pc23[33]);
FA1A GS23_34(ps24[33], pc24[34], g23[34], ps23[34], pc23[34]);
FA1A GS23_35(ps24[34], pc24[35], g23[35], ps23[35], pc23[35]);
FA1A GS23_36(ps24[35], pc24[36], g23[36], ps23[36], pc23[36]);
FA1A GS23_37(ps24[36], pc24[37], g23[37], ps23[37], pc23[37]);
FA1A GS23_38(ps24[37], pc24[38], g23[38], ps23[38], pc23[38]);
FA1A GS23_39(ps24[38], pc24[39], g23[39], ps23[39], pc23[39]);
FA1A GS23_40(ps24[39], pc24[40], g23[40], ps23[40], pc23[40]);
FA1A GS23_41(ps24[40], pc24[41], g23[41], ps23[41], pc23[41]);
FA1A GS23_42(ps24[41], pc24[42], g23[42], ps23[42], pc23[42]);
FA1A GS23_43(ps24[42], pc24[43], g23[43], ps23[43], pc23[43]);
FA1A GS23_44(ps24[43], pc24[44], g23[44], ps23[44], pc23[44]);
FA1A GS23_45(ps24[44], pc24[45], g23[45], ps23[45], pc23[45]);
FA1A GS23_46(ps24[45], pc24[46], g23[46], ps23[46], pc23[46]);
FA1A GS23_47(ps24[46], pc24[47], g23[47], ps23[47], pc23[47]);
FA1A GS23_48(ps24[47], pc24[48], g23[48], ps23[48], pc23[48]);
FA1A GS23_49(ps24[48], pc24[49], g23[49], ps23[49], pc23[49]);
FA1A GS23_50(ps24[49], pc24[50], g23[50], ps23[50], pc23[50]);
FA1A GS23_51(ps24[50], pc24[51], g23[51], ps23[51], pc23[51]);
FA1A GS23_52(ps24[51], pc24[52], g23[52], ps23[52], pc23[52]);
FA1A GS23_53(ps24[52], pc24[53], g23[53], ps23[53], pc23[53]);
FA1A GS23_54(ps24[53], pc24[54], g23[54], ps23[54], pc23[54]);
FA1A GS23_55(ps24[54], pc24[55], g23[55], ps23[55], pc23[55]);
FA1A GS23_56(ps24[55], pc24[56], g23[56], ps23[56], pc23[56]);
FA1A GS23_57(ps24[56], pc24[57], g23[57], ps23[57], pc23[57]);
FA1A GS23_58(ps24[57], pc24[58], g23[58], ps23[58], pc23[58]);
FA1A GS23_59(ps24[58], pc24[59], g23[59], ps23[59], pc23[59]);
FA1A GS23_60(ps24[59], pc24[60], g23[60], ps23[60], pc23[60]);
FA1A GS23_61(ps24[60], pc24[61], g23[61], ps23[61], pc23[61]);
FA1A GS23_62(ps24[61], pc24[62], g23[62], ps23[62], pc23[62]);
FA1A GS23_63(ps24[62], pc24[63], g23[63], ps23[63], pc23[63]);
FA1A GS22_9(g23[8], pc23[9], g22[9], ps22[9], pc22[9]);
FA1A GS22_10(ps23[9], pc23[10], g22[10], ps22[10], pc22[10]);
FA1A GS22_11(ps23[10], pc23[11], g22[11], ps22[11], pc22[11]);
FA1A GS22_12(ps23[11], pc23[12], g22[12], ps22[12], pc22[12]);
FA1A GS22_13(ps23[12], pc23[13], g22[13], ps22[13], pc22[13]);
FA1A GS22_14(ps23[13], pc23[14], g22[14], ps22[14], pc22[14]);
FA1A GS22_15(ps23[14], pc23[15], g22[15], ps22[15], pc22[15]);
FA1A GS22_16(ps23[15], pc23[16], g22[16], ps22[16], pc22[16]);
FA1A GS22_17(ps23[16], pc23[17], g22[17], ps22[17], pc22[17]);
FA1A GS22_18(ps23[17], pc23[18], g22[18], ps22[18], pc22[18]);
FA1A GS22_19(ps23[18], pc23[19], g22[19], ps22[19], pc22[19]);
FA1A GS22_20(ps23[19], pc23[20], g22[20], ps22[20], pc22[20]);
FA1A GS22_21(ps23[20], pc23[21], g22[21], ps22[21], pc22[21]);
FA1A GS22_22(ps23[21], pc23[22], g22[22], ps22[22], pc22[22]);
FA1A GS22_23(ps23[22], pc23[23], g22[23], ps22[23], pc22[23]);
FA1A GS22_24(ps23[23], pc23[24], g22[24], ps22[24], pc22[24]);
FA1A GS22_25(ps23[24], pc23[25], g22[25], ps22[25], pc22[25]);
FA1A GS22_26(ps23[25], pc23[26], g22[26], ps22[26], pc22[26]);
FA1A GS22_27(ps23[26], pc23[27], g22[27], ps22[27], pc22[27]);
FA1A GS22_28(ps23[27], pc23[28], g22[28], ps22[28], pc22[28]);
FA1A GS22_29(ps23[28], pc23[29], g22[29], ps22[29], pc22[29]);
FA1A GS22_30(ps23[29], pc23[30], g22[30], ps22[30], pc22[30]);
FA1A GS22_31(ps23[30], pc23[31], g22[31], ps22[31], pc22[31]);
FA1A GS22_32(ps23[31], pc23[32], g22[32], ps22[32], pc22[32]);
FA1A GS22_33(ps23[32], pc23[33], g22[33], ps22[33], pc22[33]);
FA1A GS22_34(ps23[33], pc23[34], g22[34], ps22[34], pc22[34]);
FA1A GS22_35(ps23[34], pc23[35], g22[35], ps22[35], pc22[35]);
FA1A GS22_36(ps23[35], pc23[36], g22[36], ps22[36], pc22[36]);
FA1A GS22_37(ps23[36], pc23[37], g22[37], ps22[37], pc22[37]);
FA1A GS22_38(ps23[37], pc23[38], g22[38], ps22[38], pc22[38]);
FA1A GS22_39(ps23[38], pc23[39], g22[39], ps22[39], pc22[39]);
FA1A GS22_40(ps23[39], pc23[40], g22[40], ps22[40], pc22[40]);
FA1A GS22_41(ps23[40], pc23[41], g22[41], ps22[41], pc22[41]);
FA1A GS22_42(ps23[41], pc23[42], g22[42], ps22[42], pc22[42]);
FA1A GS22_43(ps23[42], pc23[43], g22[43], ps22[43], pc22[43]);
FA1A GS22_44(ps23[43], pc23[44], g22[44], ps22[44], pc22[44]);
FA1A GS22_45(ps23[44], pc23[45], g22[45], ps22[45], pc22[45]);
FA1A GS22_46(ps23[45], pc23[46], g22[46], ps22[46], pc22[46]);
FA1A GS22_47(ps23[46], pc23[47], g22[47], ps22[47], pc22[47]);
FA1A GS22_48(ps23[47], pc23[48], g22[48], ps22[48], pc22[48]);
FA1A GS22_49(ps23[48], pc23[49], g22[49], ps22[49], pc22[49]);
FA1A GS22_50(ps23[49], pc23[50], g22[50], ps22[50], pc22[50]);
FA1A GS22_51(ps23[50], pc23[51], g22[51], ps22[51], pc22[51]);
FA1A GS22_52(ps23[51], pc23[52], g22[52], ps22[52], pc22[52]);
FA1A GS22_53(ps23[52], pc23[53], g22[53], ps22[53], pc22[53]);
FA1A GS22_54(ps23[53], pc23[54], g22[54], ps22[54], pc22[54]);
FA1A GS22_55(ps23[54], pc23[55], g22[55], ps22[55], pc22[55]);
FA1A GS22_56(ps23[55], pc23[56], g22[56], ps22[56], pc22[56]);
FA1A GS22_57(ps23[56], pc23[57], g22[57], ps22[57], pc22[57]);
FA1A GS22_58(ps23[57], pc23[58], g22[58], ps22[58], pc22[58]);
FA1A GS22_59(ps23[58], pc23[59], g22[59], ps22[59], pc22[59]);
FA1A GS22_60(ps23[59], pc23[60], g22[60], ps22[60], pc22[60]);
FA1A GS22_61(ps23[60], pc23[61], g22[61], ps22[61], pc22[61]);
FA1A GS22_62(ps23[61], pc23[62], g22[62], ps22[62], pc22[62]);
FA1A GS22_63(ps23[62], pc23[63], g22[63], ps22[63], pc22[63]);
FA1A GS21_9(g22[8], pc22[9], g21[9], ps21[9], pc21[9]);
FA1A GS21_10(ps22[9], pc22[10], g21[10], ps21[10], pc21[10]);
FA1A GS21_11(ps22[10], pc22[11], g21[11], ps21[11], pc21[11]);
FA1A GS21_12(ps22[11], pc22[12], g21[12], ps21[12], pc21[12]);
FA1A GS21_13(ps22[12], pc22[13], g21[13], ps21[13], pc21[13]);
FA1A GS21_14(ps22[13], pc22[14], g21[14], ps21[14], pc21[14]);
FA1A GS21_15(ps22[14], pc22[15], g21[15], ps21[15], pc21[15]);
FA1A GS21_16(ps22[15], pc22[16], g21[16], ps21[16], pc21[16]);
FA1A GS21_17(ps22[16], pc22[17], g21[17], ps21[17], pc21[17]);
FA1A GS21_18(ps22[17], pc22[18], g21[18], ps21[18], pc21[18]);
FA1A GS21_19(ps22[18], pc22[19], g21[19], ps21[19], pc21[19]);
FA1A GS21_20(ps22[19], pc22[20], g21[20], ps21[20], pc21[20]);
FA1A GS21_21(ps22[20], pc22[21], g21[21], ps21[21], pc21[21]);
FA1A GS21_22(ps22[21], pc22[22], g21[22], ps21[22], pc21[22]);
FA1A GS21_23(ps22[22], pc22[23], g21[23], ps21[23], pc21[23]);
FA1A GS21_24(ps22[23], pc22[24], g21[24], ps21[24], pc21[24]);
FA1A GS21_25(ps22[24], pc22[25], g21[25], ps21[25], pc21[25]);
FA1A GS21_26(ps22[25], pc22[26], g21[26], ps21[26], pc21[26]);
FA1A GS21_27(ps22[26], pc22[27], g21[27], ps21[27], pc21[27]);
FA1A GS21_28(ps22[27], pc22[28], g21[28], ps21[28], pc21[28]);
FA1A GS21_29(ps22[28], pc22[29], g21[29], ps21[29], pc21[29]);
FA1A GS21_30(ps22[29], pc22[30], g21[30], ps21[30], pc21[30]);
FA1A GS21_31(ps22[30], pc22[31], g21[31], ps21[31], pc21[31]);
FA1A GS21_32(ps22[31], pc22[32], g21[32], ps21[32], pc21[32]);
FA1A GS21_33(ps22[32], pc22[33], g21[33], ps21[33], pc21[33]);
FA1A GS21_34(ps22[33], pc22[34], g21[34], ps21[34], pc21[34]);
FA1A GS21_35(ps22[34], pc22[35], g21[35], ps21[35], pc21[35]);
FA1A GS21_36(ps22[35], pc22[36], g21[36], ps21[36], pc21[36]);
FA1A GS21_37(ps22[36], pc22[37], g21[37], ps21[37], pc21[37]);
FA1A GS21_38(ps22[37], pc22[38], g21[38], ps21[38], pc21[38]);
FA1A GS21_39(ps22[38], pc22[39], g21[39], ps21[39], pc21[39]);
FA1A GS21_40(ps22[39], pc22[40], g21[40], ps21[40], pc21[40]);
FA1A GS21_41(ps22[40], pc22[41], g21[41], ps21[41], pc21[41]);
FA1A GS21_42(ps22[41], pc22[42], g21[42], ps21[42], pc21[42]);
FA1A GS21_43(ps22[42], pc22[43], g21[43], ps21[43], pc21[43]);
FA1A GS21_44(ps22[43], pc22[44], g21[44], ps21[44], pc21[44]);
FA1A GS21_45(ps22[44], pc22[45], g21[45], ps21[45], pc21[45]);
FA1A GS21_46(ps22[45], pc22[46], g21[46], ps21[46], pc21[46]);
FA1A GS21_47(ps22[46], pc22[47], g21[47], ps21[47], pc21[47]);
FA1A GS21_48(ps22[47], pc22[48], g21[48], ps21[48], pc21[48]);
FA1A GS21_49(ps22[48], pc22[49], g21[49], ps21[49], pc21[49]);
FA1A GS21_50(ps22[49], pc22[50], g21[50], ps21[50], pc21[50]);
FA1A GS21_51(ps22[50], pc22[51], g21[51], ps21[51], pc21[51]);
FA1A GS21_52(ps22[51], pc22[52], g21[52], ps21[52], pc21[52]);
FA1A GS21_53(ps22[52], pc22[53], g21[53], ps21[53], pc21[53]);
FA1A GS21_54(ps22[53], pc22[54], g21[54], ps21[54], pc21[54]);
FA1A GS21_55(ps22[54], pc22[55], g21[55], ps21[55], pc21[55]);
FA1A GS21_56(ps22[55], pc22[56], g21[56], ps21[56], pc21[56]);
FA1A GS21_57(ps22[56], pc22[57], g21[57], ps21[57], pc21[57]);
FA1A GS21_58(ps22[57], pc22[58], g21[58], ps21[58], pc21[58]);
FA1A GS21_59(ps22[58], pc22[59], g21[59], ps21[59], pc21[59]);
FA1A GS21_60(ps22[59], pc22[60], g21[60], ps21[60], pc21[60]);
FA1A GS21_61(ps22[60], pc22[61], g21[61], ps21[61], pc21[61]);
FA1A GS21_62(ps22[61], pc22[62], g21[62], ps21[62], pc21[62]);
FA1A GS21_63(ps22[62], pc22[63], g21[63], ps21[63], pc21[63]);
FA1A GS20_9(g21[8], pc21[9], g20[9], ps20[9], pc20[9]);
FA1A GS20_10(ps21[9], pc21[10], g20[10], ps20[10], pc20[10]);
FA1A GS20_11(ps21[10], pc21[11], g20[11], ps20[11], pc20[11]);
FA1A GS20_12(ps21[11], pc21[12], g20[12], ps20[12], pc20[12]);
FA1A GS20_13(ps21[12], pc21[13], g20[13], ps20[13], pc20[13]);
FA1A GS20_14(ps21[13], pc21[14], g20[14], ps20[14], pc20[14]);
FA1A GS20_15(ps21[14], pc21[15], g20[15], ps20[15], pc20[15]);
FA1A GS20_16(ps21[15], pc21[16], g20[16], ps20[16], pc20[16]);
FA1A GS20_17(ps21[16], pc21[17], g20[17], ps20[17], pc20[17]);
FA1A GS20_18(ps21[17], pc21[18], g20[18], ps20[18], pc20[18]);
FA1A GS20_19(ps21[18], pc21[19], g20[19], ps20[19], pc20[19]);
FA1A GS20_20(ps21[19], pc21[20], g20[20], ps20[20], pc20[20]);
FA1A GS20_21(ps21[20], pc21[21], g20[21], ps20[21], pc20[21]);
FA1A GS20_22(ps21[21], pc21[22], g20[22], ps20[22], pc20[22]);
FA1A GS20_23(ps21[22], pc21[23], g20[23], ps20[23], pc20[23]);
FA1A GS20_24(ps21[23], pc21[24], g20[24], ps20[24], pc20[24]);
FA1A GS20_25(ps21[24], pc21[25], g20[25], ps20[25], pc20[25]);
FA1A GS20_26(ps21[25], pc21[26], g20[26], ps20[26], pc20[26]);
FA1A GS20_27(ps21[26], pc21[27], g20[27], ps20[27], pc20[27]);
FA1A GS20_28(ps21[27], pc21[28], g20[28], ps20[28], pc20[28]);
FA1A GS20_29(ps21[28], pc21[29], g20[29], ps20[29], pc20[29]);
FA1A GS20_30(ps21[29], pc21[30], g20[30], ps20[30], pc20[30]);
FA1A GS20_31(ps21[30], pc21[31], g20[31], ps20[31], pc20[31]);
FA1A GS20_32(ps21[31], pc21[32], g20[32], ps20[32], pc20[32]);
FA1A GS20_33(ps21[32], pc21[33], g20[33], ps20[33], pc20[33]);
FA1A GS20_34(ps21[33], pc21[34], g20[34], ps20[34], pc20[34]);
FA1A GS20_35(ps21[34], pc21[35], g20[35], ps20[35], pc20[35]);
FA1A GS20_36(ps21[35], pc21[36], g20[36], ps20[36], pc20[36]);
FA1A GS20_37(ps21[36], pc21[37], g20[37], ps20[37], pc20[37]);
FA1A GS20_38(ps21[37], pc21[38], g20[38], ps20[38], pc20[38]);
FA1A GS20_39(ps21[38], pc21[39], g20[39], ps20[39], pc20[39]);
FA1A GS20_40(ps21[39], pc21[40], g20[40], ps20[40], pc20[40]);
FA1A GS20_41(ps21[40], pc21[41], g20[41], ps20[41], pc20[41]);
FA1A GS20_42(ps21[41], pc21[42], g20[42], ps20[42], pc20[42]);
FA1A GS20_43(ps21[42], pc21[43], g20[43], ps20[43], pc20[43]);
FA1A GS20_44(ps21[43], pc21[44], g20[44], ps20[44], pc20[44]);
FA1A GS20_45(ps21[44], pc21[45], g20[45], ps20[45], pc20[45]);
FA1A GS20_46(ps21[45], pc21[46], g20[46], ps20[46], pc20[46]);
FA1A GS20_47(ps21[46], pc21[47], g20[47], ps20[47], pc20[47]);
FA1A GS20_48(ps21[47], pc21[48], g20[48], ps20[48], pc20[48]);
FA1A GS20_49(ps21[48], pc21[49], g20[49], ps20[49], pc20[49]);
FA1A GS20_50(ps21[49], pc21[50], g20[50], ps20[50], pc20[50]);
FA1A GS20_51(ps21[50], pc21[51], g20[51], ps20[51], pc20[51]);
FA1A GS20_52(ps21[51], pc21[52], g20[52], ps20[52], pc20[52]);
FA1A GS20_53(ps21[52], pc21[53], g20[53], ps20[53], pc20[53]);
FA1A GS20_54(ps21[53], pc21[54], g20[54], ps20[54], pc20[54]);
FA1A GS20_55(ps21[54], pc21[55], g20[55], ps20[55], pc20[55]);
FA1A GS20_56(ps21[55], pc21[56], g20[56], ps20[56], pc20[56]);
FA1A GS20_57(ps21[56], pc21[57], g20[57], ps20[57], pc20[57]);
FA1A GS20_58(ps21[57], pc21[58], g20[58], ps20[58], pc20[58]);
FA1A GS20_59(ps21[58], pc21[59], g20[59], ps20[59], pc20[59]);
FA1A GS20_60(ps21[59], pc21[60], g20[60], ps20[60], pc20[60]);
FA1A GS20_61(ps21[60], pc21[61], g20[61], ps20[61], pc20[61]);
FA1A GS20_62(ps21[61], pc21[62], g20[62], ps20[62], pc20[62]);
FA1A GS20_63(ps21[62], pc21[63], g20[63], ps20[63], pc20[63]);
FA1A GS19_9(g20[8], pc20[9], g19[9], ps19[9], pc19[9]);
FA1A GS19_10(ps20[9], pc20[10], g19[10], ps19[10], pc19[10]);
FA1A GS19_11(ps20[10], pc20[11], g19[11], ps19[11], pc19[11]);
FA1A GS19_12(ps20[11], pc20[12], g19[12], ps19[12], pc19[12]);
FA1A GS19_13(ps20[12], pc20[13], g19[13], ps19[13], pc19[13]);
FA1A GS19_14(ps20[13], pc20[14], g19[14], ps19[14], pc19[14]);
FA1A GS19_15(ps20[14], pc20[15], g19[15], ps19[15], pc19[15]);
FA1A GS19_16(ps20[15], pc20[16], g19[16], ps19[16], pc19[16]);
FA1A GS19_17(ps20[16], pc20[17], g19[17], ps19[17], pc19[17]);
FA1A GS19_18(ps20[17], pc20[18], g19[18], ps19[18], pc19[18]);
FA1A GS19_19(ps20[18], pc20[19], g19[19], ps19[19], pc19[19]);
FA1A GS19_20(ps20[19], pc20[20], g19[20], ps19[20], pc19[20]);
FA1A GS19_21(ps20[20], pc20[21], g19[21], ps19[21], pc19[21]);
FA1A GS19_22(ps20[21], pc20[22], g19[22], ps19[22], pc19[22]);
FA1A GS19_23(ps20[22], pc20[23], g19[23], ps19[23], pc19[23]);
FA1A GS19_24(ps20[23], pc20[24], g19[24], ps19[24], pc19[24]);
FA1A GS19_25(ps20[24], pc20[25], g19[25], ps19[25], pc19[25]);
FA1A GS19_26(ps20[25], pc20[26], g19[26], ps19[26], pc19[26]);
FA1A GS19_27(ps20[26], pc20[27], g19[27], ps19[27], pc19[27]);
FA1A GS19_28(ps20[27], pc20[28], g19[28], ps19[28], pc19[28]);
FA1A GS19_29(ps20[28], pc20[29], g19[29], ps19[29], pc19[29]);
FA1A GS19_30(ps20[29], pc20[30], g19[30], ps19[30], pc19[30]);
FA1A GS19_31(ps20[30], pc20[31], g19[31], ps19[31], pc19[31]);
FA1A GS19_32(ps20[31], pc20[32], g19[32], ps19[32], pc19[32]);
FA1A GS19_33(ps20[32], pc20[33], g19[33], ps19[33], pc19[33]);
FA1A GS19_34(ps20[33], pc20[34], g19[34], ps19[34], pc19[34]);
FA1A GS19_35(ps20[34], pc20[35], g19[35], ps19[35], pc19[35]);
FA1A GS19_36(ps20[35], pc20[36], g19[36], ps19[36], pc19[36]);
FA1A GS19_37(ps20[36], pc20[37], g19[37], ps19[37], pc19[37]);
FA1A GS19_38(ps20[37], pc20[38], g19[38], ps19[38], pc19[38]);
FA1A GS19_39(ps20[38], pc20[39], g19[39], ps19[39], pc19[39]);
FA1A GS19_40(ps20[39], pc20[40], g19[40], ps19[40], pc19[40]);
FA1A GS19_41(ps20[40], pc20[41], g19[41], ps19[41], pc19[41]);
FA1A GS19_42(ps20[41], pc20[42], g19[42], ps19[42], pc19[42]);
FA1A GS19_43(ps20[42], pc20[43], g19[43], ps19[43], pc19[43]);
FA1A GS19_44(ps20[43], pc20[44], g19[44], ps19[44], pc19[44]);
FA1A GS19_45(ps20[44], pc20[45], g19[45], ps19[45], pc19[45]);
FA1A GS19_46(ps20[45], pc20[46], g19[46], ps19[46], pc19[46]);
FA1A GS19_47(ps20[46], pc20[47], g19[47], ps19[47], pc19[47]);
FA1A GS19_48(ps20[47], pc20[48], g19[48], ps19[48], pc19[48]);
FA1A GS19_49(ps20[48], pc20[49], g19[49], ps19[49], pc19[49]);
FA1A GS19_50(ps20[49], pc20[50], g19[50], ps19[50], pc19[50]);
FA1A GS19_51(ps20[50], pc20[51], g19[51], ps19[51], pc19[51]);
FA1A GS19_52(ps20[51], pc20[52], g19[52], ps19[52], pc19[52]);
FA1A GS19_53(ps20[52], pc20[53], g19[53], ps19[53], pc19[53]);
FA1A GS19_54(ps20[53], pc20[54], g19[54], ps19[54], pc19[54]);
FA1A GS19_55(ps20[54], pc20[55], g19[55], ps19[55], pc19[55]);
FA1A GS19_56(ps20[55], pc20[56], g19[56], ps19[56], pc19[56]);
FA1A GS19_57(ps20[56], pc20[57], g19[57], ps19[57], pc19[57]);
FA1A GS19_58(ps20[57], pc20[58], g19[58], ps19[58], pc19[58]);
FA1A GS19_59(ps20[58], pc20[59], g19[59], ps19[59], pc19[59]);
FA1A GS19_60(ps20[59], pc20[60], g19[60], ps19[60], pc19[60]);
FA1A GS19_61(ps20[60], pc20[61], g19[61], ps19[61], pc19[61]);
FA1A GS19_62(ps20[61], pc20[62], g19[62], ps19[62], pc19[62]);
FA1A GS19_63(ps20[62], pc20[63], g19[63], ps19[63], pc19[63]);
FA1A GS18_9(g19[8], pc19[9], g18[9], ps18[9], pc18[9]);
FA1A GS18_10(ps19[9], pc19[10], g18[10], ps18[10], pc18[10]);
FA1A GS18_11(ps19[10], pc19[11], g18[11], ps18[11], pc18[11]);
FA1A GS18_12(ps19[11], pc19[12], g18[12], ps18[12], pc18[12]);
FA1A GS18_13(ps19[12], pc19[13], g18[13], ps18[13], pc18[13]);
FA1A GS18_14(ps19[13], pc19[14], g18[14], ps18[14], pc18[14]);
FA1A GS18_15(ps19[14], pc19[15], g18[15], ps18[15], pc18[15]);
FA1A GS18_16(ps19[15], pc19[16], g18[16], ps18[16], pc18[16]);
FA1A GS18_17(ps19[16], pc19[17], g18[17], ps18[17], pc18[17]);
FA1A GS18_18(ps19[17], pc19[18], g18[18], ps18[18], pc18[18]);
FA1A GS18_19(ps19[18], pc19[19], g18[19], ps18[19], pc18[19]);
FA1A GS18_20(ps19[19], pc19[20], g18[20], ps18[20], pc18[20]);
FA1A GS18_21(ps19[20], pc19[21], g18[21], ps18[21], pc18[21]);
FA1A GS18_22(ps19[21], pc19[22], g18[22], ps18[22], pc18[22]);
FA1A GS18_23(ps19[22], pc19[23], g18[23], ps18[23], pc18[23]);
FA1A GS18_24(ps19[23], pc19[24], g18[24], ps18[24], pc18[24]);
FA1A GS18_25(ps19[24], pc19[25], g18[25], ps18[25], pc18[25]);
FA1A GS18_26(ps19[25], pc19[26], g18[26], ps18[26], pc18[26]);
FA1A GS18_27(ps19[26], pc19[27], g18[27], ps18[27], pc18[27]);
FA1A GS18_28(ps19[27], pc19[28], g18[28], ps18[28], pc18[28]);
FA1A GS18_29(ps19[28], pc19[29], g18[29], ps18[29], pc18[29]);
FA1A GS18_30(ps19[29], pc19[30], g18[30], ps18[30], pc18[30]);
FA1A GS18_31(ps19[30], pc19[31], g18[31], ps18[31], pc18[31]);
FA1A GS18_32(ps19[31], pc19[32], g18[32], ps18[32], pc18[32]);
FA1A GS18_33(ps19[32], pc19[33], g18[33], ps18[33], pc18[33]);
FA1A GS18_34(ps19[33], pc19[34], g18[34], ps18[34], pc18[34]);
FA1A GS18_35(ps19[34], pc19[35], g18[35], ps18[35], pc18[35]);
FA1A GS18_36(ps19[35], pc19[36], g18[36], ps18[36], pc18[36]);
FA1A GS18_37(ps19[36], pc19[37], g18[37], ps18[37], pc18[37]);
FA1A GS18_38(ps19[37], pc19[38], g18[38], ps18[38], pc18[38]);
FA1A GS18_39(ps19[38], pc19[39], g18[39], ps18[39], pc18[39]);
FA1A GS18_40(ps19[39], pc19[40], g18[40], ps18[40], pc18[40]);
FA1A GS18_41(ps19[40], pc19[41], g18[41], ps18[41], pc18[41]);
FA1A GS18_42(ps19[41], pc19[42], g18[42], ps18[42], pc18[42]);
FA1A GS18_43(ps19[42], pc19[43], g18[43], ps18[43], pc18[43]);
FA1A GS18_44(ps19[43], pc19[44], g18[44], ps18[44], pc18[44]);
FA1A GS18_45(ps19[44], pc19[45], g18[45], ps18[45], pc18[45]);
FA1A GS18_46(ps19[45], pc19[46], g18[46], ps18[46], pc18[46]);
FA1A GS18_47(ps19[46], pc19[47], g18[47], ps18[47], pc18[47]);
FA1A GS18_48(ps19[47], pc19[48], g18[48], ps18[48], pc18[48]);
FA1A GS18_49(ps19[48], pc19[49], g18[49], ps18[49], pc18[49]);
FA1A GS18_50(ps19[49], pc19[50], g18[50], ps18[50], pc18[50]);
FA1A GS18_51(ps19[50], pc19[51], g18[51], ps18[51], pc18[51]);
FA1A GS18_52(ps19[51], pc19[52], g18[52], ps18[52], pc18[52]);
FA1A GS18_53(ps19[52], pc19[53], g18[53], ps18[53], pc18[53]);
FA1A GS18_54(ps19[53], pc19[54], g18[54], ps18[54], pc18[54]);
FA1A GS18_55(ps19[54], pc19[55], g18[55], ps18[55], pc18[55]);
FA1A GS18_56(ps19[55], pc19[56], g18[56], ps18[56], pc18[56]);
FA1A GS18_57(ps19[56], pc19[57], g18[57], ps18[57], pc18[57]);
FA1A GS18_58(ps19[57], pc19[58], g18[58], ps18[58], pc18[58]);
FA1A GS18_59(ps19[58], pc19[59], g18[59], ps18[59], pc18[59]);
FA1A GS18_60(ps19[59], pc19[60], g18[60], ps18[60], pc18[60]);
FA1A GS18_61(ps19[60], pc19[61], g18[61], ps18[61], pc18[61]);
FA1A GS18_62(ps19[61], pc19[62], g18[62], ps18[62], pc18[62]);
FA1A GS18_63(ps19[62], pc19[63], g18[63], ps18[63], pc18[63]);
FA1A GS17_9(g18[8], pc18[9], g17[9], ps17[9], pc17[9]);
FA1A GS17_10(ps18[9], pc18[10], g17[10], ps17[10], pc17[10]);
FA1A GS17_11(ps18[10], pc18[11], g17[11], ps17[11], pc17[11]);
FA1A GS17_12(ps18[11], pc18[12], g17[12], ps17[12], pc17[12]);
FA1A GS17_13(ps18[12], pc18[13], g17[13], ps17[13], pc17[13]);
FA1A GS17_14(ps18[13], pc18[14], g17[14], ps17[14], pc17[14]);
FA1A GS17_15(ps18[14], pc18[15], g17[15], ps17[15], pc17[15]);
FA1A GS17_16(ps18[15], pc18[16], g17[16], ps17[16], pc17[16]);
FA1A GS17_17(ps18[16], pc18[17], g17[17], ps17[17], pc17[17]);
FA1A GS17_18(ps18[17], pc18[18], g17[18], ps17[18], pc17[18]);
FA1A GS17_19(ps18[18], pc18[19], g17[19], ps17[19], pc17[19]);
FA1A GS17_20(ps18[19], pc18[20], g17[20], ps17[20], pc17[20]);
FA1A GS17_21(ps18[20], pc18[21], g17[21], ps17[21], pc17[21]);
FA1A GS17_22(ps18[21], pc18[22], g17[22], ps17[22], pc17[22]);
FA1A GS17_23(ps18[22], pc18[23], g17[23], ps17[23], pc17[23]);
FA1A GS17_24(ps18[23], pc18[24], g17[24], ps17[24], pc17[24]);
FA1A GS17_25(ps18[24], pc18[25], g17[25], ps17[25], pc17[25]);
FA1A GS17_26(ps18[25], pc18[26], g17[26], ps17[26], pc17[26]);
FA1A GS17_27(ps18[26], pc18[27], g17[27], ps17[27], pc17[27]);
FA1A GS17_28(ps18[27], pc18[28], g17[28], ps17[28], pc17[28]);
FA1A GS17_29(ps18[28], pc18[29], g17[29], ps17[29], pc17[29]);
FA1A GS17_30(ps18[29], pc18[30], g17[30], ps17[30], pc17[30]);
FA1A GS17_31(ps18[30], pc18[31], g17[31], ps17[31], pc17[31]);
FA1A GS17_32(ps18[31], pc18[32], g17[32], ps17[32], pc17[32]);
FA1A GS17_33(ps18[32], pc18[33], g17[33], ps17[33], pc17[33]);
FA1A GS17_34(ps18[33], pc18[34], g17[34], ps17[34], pc17[34]);
FA1A GS17_35(ps18[34], pc18[35], g17[35], ps17[35], pc17[35]);
FA1A GS17_36(ps18[35], pc18[36], g17[36], ps17[36], pc17[36]);
FA1A GS17_37(ps18[36], pc18[37], g17[37], ps17[37], pc17[37]);
FA1A GS17_38(ps18[37], pc18[38], g17[38], ps17[38], pc17[38]);
FA1A GS17_39(ps18[38], pc18[39], g17[39], ps17[39], pc17[39]);
FA1A GS17_40(ps18[39], pc18[40], g17[40], ps17[40], pc17[40]);
FA1A GS17_41(ps18[40], pc18[41], g17[41], ps17[41], pc17[41]);
FA1A GS17_42(ps18[41], pc18[42], g17[42], ps17[42], pc17[42]);
FA1A GS17_43(ps18[42], pc18[43], g17[43], ps17[43], pc17[43]);
FA1A GS17_44(ps18[43], pc18[44], g17[44], ps17[44], pc17[44]);
FA1A GS17_45(ps18[44], pc18[45], g17[45], ps17[45], pc17[45]);
FA1A GS17_46(ps18[45], pc18[46], g17[46], ps17[46], pc17[46]);
FA1A GS17_47(ps18[46], pc18[47], g17[47], ps17[47], pc17[47]);
FA1A GS17_48(ps18[47], pc18[48], g17[48], ps17[48], pc17[48]);
FA1A GS17_49(ps18[48], pc18[49], g17[49], ps17[49], pc17[49]);
FA1A GS17_50(ps18[49], pc18[50], g17[50], ps17[50], pc17[50]);
FA1A GS17_51(ps18[50], pc18[51], g17[51], ps17[51], pc17[51]);
FA1A GS17_52(ps18[51], pc18[52], g17[52], ps17[52], pc17[52]);
FA1A GS17_53(ps18[52], pc18[53], g17[53], ps17[53], pc17[53]);
FA1A GS17_54(ps18[53], pc18[54], g17[54], ps17[54], pc17[54]);
FA1A GS17_55(ps18[54], pc18[55], g17[55], ps17[55], pc17[55]);
FA1A GS17_56(ps18[55], pc18[56], g17[56], ps17[56], pc17[56]);
FA1A GS17_57(ps18[56], pc18[57], g17[57], ps17[57], pc17[57]);
FA1A GS17_58(ps18[57], pc18[58], g17[58], ps17[58], pc17[58]);
FA1A GS17_59(ps18[58], pc18[59], g17[59], ps17[59], pc17[59]);
FA1A GS17_60(ps18[59], pc18[60], g17[60], ps17[60], pc17[60]);
FA1A GS17_61(ps18[60], pc18[61], g17[61], ps17[61], pc17[61]);
FA1A GS17_62(ps18[61], pc18[62], g17[62], ps17[62], pc17[62]);
FA1A GS17_63(ps18[62], pc18[63], g17[63], ps17[63], pc17[63]);
FA1A GS16_9(g17[8], pc17[9], g16[9], ps16[9], pc16[9]);
FA1A GS16_10(ps17[9], pc17[10], g16[10], ps16[10], pc16[10]);
FA1A GS16_11(ps17[10], pc17[11], g16[11], ps16[11], pc16[11]);
FA1A GS16_12(ps17[11], pc17[12], g16[12], ps16[12], pc16[12]);
FA1A GS16_13(ps17[12], pc17[13], g16[13], ps16[13], pc16[13]);
FA1A GS16_14(ps17[13], pc17[14], g16[14], ps16[14], pc16[14]);
FA1A GS16_15(ps17[14], pc17[15], g16[15], ps16[15], pc16[15]);
FA1A GS16_16(ps17[15], pc17[16], g16[16], ps16[16], pc16[16]);
FA1A GS16_17(ps17[16], pc17[17], g16[17], ps16[17], pc16[17]);
FA1A GS16_18(ps17[17], pc17[18], g16[18], ps16[18], pc16[18]);
FA1A GS16_19(ps17[18], pc17[19], g16[19], ps16[19], pc16[19]);
FA1A GS16_20(ps17[19], pc17[20], g16[20], ps16[20], pc16[20]);
FA1A GS16_21(ps17[20], pc17[21], g16[21], ps16[21], pc16[21]);
FA1A GS16_22(ps17[21], pc17[22], g16[22], ps16[22], pc16[22]);
FA1A GS16_23(ps17[22], pc17[23], g16[23], ps16[23], pc16[23]);
FA1A GS16_24(ps17[23], pc17[24], g16[24], ps16[24], pc16[24]);
FA1A GS16_25(ps17[24], pc17[25], g16[25], ps16[25], pc16[25]);
FA1A GS16_26(ps17[25], pc17[26], g16[26], ps16[26], pc16[26]);
FA1A GS16_27(ps17[26], pc17[27], g16[27], ps16[27], pc16[27]);
FA1A GS16_28(ps17[27], pc17[28], g16[28], ps16[28], pc16[28]);
FA1A GS16_29(ps17[28], pc17[29], g16[29], ps16[29], pc16[29]);
FA1A GS16_30(ps17[29], pc17[30], g16[30], ps16[30], pc16[30]);
FA1A GS16_31(ps17[30], pc17[31], g16[31], ps16[31], pc16[31]);
FA1A GS16_32(ps17[31], pc17[32], g16[32], ps16[32], pc16[32]);
FA1A GS16_33(ps17[32], pc17[33], g16[33], ps16[33], pc16[33]);
FA1A GS16_34(ps17[33], pc17[34], g16[34], ps16[34], pc16[34]);
FA1A GS16_35(ps17[34], pc17[35], g16[35], ps16[35], pc16[35]);
FA1A GS16_36(ps17[35], pc17[36], g16[36], ps16[36], pc16[36]);
FA1A GS16_37(ps17[36], pc17[37], g16[37], ps16[37], pc16[37]);
FA1A GS16_38(ps17[37], pc17[38], g16[38], ps16[38], pc16[38]);
FA1A GS16_39(ps17[38], pc17[39], g16[39], ps16[39], pc16[39]);
FA1A GS16_40(ps17[39], pc17[40], g16[40], ps16[40], pc16[40]);
FA1A GS16_41(ps17[40], pc17[41], g16[41], ps16[41], pc16[41]);
FA1A GS16_42(ps17[41], pc17[42], g16[42], ps16[42], pc16[42]);
FA1A GS16_43(ps17[42], pc17[43], g16[43], ps16[43], pc16[43]);
FA1A GS16_44(ps17[43], pc17[44], g16[44], ps16[44], pc16[44]);
FA1A GS16_45(ps17[44], pc17[45], g16[45], ps16[45], pc16[45]);
FA1A GS16_46(ps17[45], pc17[46], g16[46], ps16[46], pc16[46]);
FA1A GS16_47(ps17[46], pc17[47], g16[47], ps16[47], pc16[47]);
FA1A GS16_48(ps17[47], pc17[48], g16[48], ps16[48], pc16[48]);
FA1A GS16_49(ps17[48], pc17[49], g16[49], ps16[49], pc16[49]);
FA1A GS16_50(ps17[49], pc17[50], g16[50], ps16[50], pc16[50]);
FA1A GS16_51(ps17[50], pc17[51], g16[51], ps16[51], pc16[51]);
FA1A GS16_52(ps17[51], pc17[52], g16[52], ps16[52], pc16[52]);
FA1A GS16_53(ps17[52], pc17[53], g16[53], ps16[53], pc16[53]);
FA1A GS16_54(ps17[53], pc17[54], g16[54], ps16[54], pc16[54]);
FA1A GS16_55(ps17[54], pc17[55], g16[55], ps16[55], pc16[55]);
FA1A GS16_56(ps17[55], pc17[56], g16[56], ps16[56], pc16[56]);
FA1A GS16_57(ps17[56], pc17[57], g16[57], ps16[57], pc16[57]);
FA1A GS16_58(ps17[57], pc17[58], g16[58], ps16[58], pc16[58]);
FA1A GS16_59(ps17[58], pc17[59], g16[59], ps16[59], pc16[59]);
FA1A GS16_60(ps17[59], pc17[60], g16[60], ps16[60], pc16[60]);
FA1A GS16_61(ps17[60], pc17[61], g16[61], ps16[61], pc16[61]);
FA1A GS16_62(ps17[61], pc17[62], g16[62], ps16[62], pc16[62]);
FA1A GS16_63(ps17[62], pc17[63], g16[63], ps16[63], pc16[63]);
FA1A GS15_9(g16[8], pc16[9], g15[9], ps15[9], pc15[9]);
FA1A GS15_10(ps16[9], pc16[10], g15[10], ps15[10], pc15[10]);
FA1A GS15_11(ps16[10], pc16[11], g15[11], ps15[11], pc15[11]);
FA1A GS15_12(ps16[11], pc16[12], g15[12], ps15[12], pc15[12]);
FA1A GS15_13(ps16[12], pc16[13], g15[13], ps15[13], pc15[13]);
FA1A GS15_14(ps16[13], pc16[14], g15[14], ps15[14], pc15[14]);
FA1A GS15_15(ps16[14], pc16[15], g15[15], ps15[15], pc15[15]);
FA1A GS15_16(ps16[15], pc16[16], g15[16], ps15[16], pc15[16]);
FA1A GS15_17(ps16[16], pc16[17], g15[17], ps15[17], pc15[17]);
FA1A GS15_18(ps16[17], pc16[18], g15[18], ps15[18], pc15[18]);
FA1A GS15_19(ps16[18], pc16[19], g15[19], ps15[19], pc15[19]);
FA1A GS15_20(ps16[19], pc16[20], g15[20], ps15[20], pc15[20]);
FA1A GS15_21(ps16[20], pc16[21], g15[21], ps15[21], pc15[21]);
FA1A GS15_22(ps16[21], pc16[22], g15[22], ps15[22], pc15[22]);
FA1A GS15_23(ps16[22], pc16[23], g15[23], ps15[23], pc15[23]);
FA1A GS15_24(ps16[23], pc16[24], g15[24], ps15[24], pc15[24]);
FA1A GS15_25(ps16[24], pc16[25], g15[25], ps15[25], pc15[25]);
FA1A GS15_26(ps16[25], pc16[26], g15[26], ps15[26], pc15[26]);
FA1A GS15_27(ps16[26], pc16[27], g15[27], ps15[27], pc15[27]);
FA1A GS15_28(ps16[27], pc16[28], g15[28], ps15[28], pc15[28]);
FA1A GS15_29(ps16[28], pc16[29], g15[29], ps15[29], pc15[29]);
FA1A GS15_30(ps16[29], pc16[30], g15[30], ps15[30], pc15[30]);
FA1A GS15_31(ps16[30], pc16[31], g15[31], ps15[31], pc15[31]);
FA1A GS15_32(ps16[31], pc16[32], g15[32], ps15[32], pc15[32]);
FA1A GS15_33(ps16[32], pc16[33], g15[33], ps15[33], pc15[33]);
FA1A GS15_34(ps16[33], pc16[34], g15[34], ps15[34], pc15[34]);
FA1A GS15_35(ps16[34], pc16[35], g15[35], ps15[35], pc15[35]);
FA1A GS15_36(ps16[35], pc16[36], g15[36], ps15[36], pc15[36]);
FA1A GS15_37(ps16[36], pc16[37], g15[37], ps15[37], pc15[37]);
FA1A GS15_38(ps16[37], pc16[38], g15[38], ps15[38], pc15[38]);
FA1A GS15_39(ps16[38], pc16[39], g15[39], ps15[39], pc15[39]);
FA1A GS15_40(ps16[39], pc16[40], g15[40], ps15[40], pc15[40]);
FA1A GS15_41(ps16[40], pc16[41], g15[41], ps15[41], pc15[41]);
FA1A GS15_42(ps16[41], pc16[42], g15[42], ps15[42], pc15[42]);
FA1A GS15_43(ps16[42], pc16[43], g15[43], ps15[43], pc15[43]);
FA1A GS15_44(ps16[43], pc16[44], g15[44], ps15[44], pc15[44]);
FA1A GS15_45(ps16[44], pc16[45], g15[45], ps15[45], pc15[45]);
FA1A GS15_46(ps16[45], pc16[46], g15[46], ps15[46], pc15[46]);
FA1A GS15_47(ps16[46], pc16[47], g15[47], ps15[47], pc15[47]);
FA1A GS15_48(ps16[47], pc16[48], g15[48], ps15[48], pc15[48]);
FA1A GS15_49(ps16[48], pc16[49], g15[49], ps15[49], pc15[49]);
FA1A GS15_50(ps16[49], pc16[50], g15[50], ps15[50], pc15[50]);
FA1A GS15_51(ps16[50], pc16[51], g15[51], ps15[51], pc15[51]);
FA1A GS15_52(ps16[51], pc16[52], g15[52], ps15[52], pc15[52]);
FA1A GS15_53(ps16[52], pc16[53], g15[53], ps15[53], pc15[53]);
FA1A GS15_54(ps16[53], pc16[54], g15[54], ps15[54], pc15[54]);
FA1A GS15_55(ps16[54], pc16[55], g15[55], ps15[55], pc15[55]);
FA1A GS15_56(ps16[55], pc16[56], g15[56], ps15[56], pc15[56]);
FA1A GS15_57(ps16[56], pc16[57], g15[57], ps15[57], pc15[57]);
FA1A GS15_58(ps16[57], pc16[58], g15[58], ps15[58], pc15[58]);
FA1A GS15_59(ps16[58], pc16[59], g15[59], ps15[59], pc15[59]);
FA1A GS15_60(ps16[59], pc16[60], g15[60], ps15[60], pc15[60]);
FA1A GS15_61(ps16[60], pc16[61], g15[61], ps15[61], pc15[61]);
FA1A GS15_62(ps16[61], pc16[62], g15[62], ps15[62], pc15[62]);
FA1A GS15_63(ps16[62], pc16[63], g15[63], ps15[63], pc15[63]);
FA1A GS14_9(g15[8], pc15[9], g14[9], ps14[9], pc14[9]);
FA1A GS14_10(ps15[9], pc15[10], g14[10], ps14[10], pc14[10]);
FA1A GS14_11(ps15[10], pc15[11], g14[11], ps14[11], pc14[11]);
FA1A GS14_12(ps15[11], pc15[12], g14[12], ps14[12], pc14[12]);
FA1A GS14_13(ps15[12], pc15[13], g14[13], ps14[13], pc14[13]);
FA1A GS14_14(ps15[13], pc15[14], g14[14], ps14[14], pc14[14]);
FA1A GS14_15(ps15[14], pc15[15], g14[15], ps14[15], pc14[15]);
FA1A GS14_16(ps15[15], pc15[16], g14[16], ps14[16], pc14[16]);
FA1A GS14_17(ps15[16], pc15[17], g14[17], ps14[17], pc14[17]);
FA1A GS14_18(ps15[17], pc15[18], g14[18], ps14[18], pc14[18]);
FA1A GS14_19(ps15[18], pc15[19], g14[19], ps14[19], pc14[19]);
FA1A GS14_20(ps15[19], pc15[20], g14[20], ps14[20], pc14[20]);
FA1A GS14_21(ps15[20], pc15[21], g14[21], ps14[21], pc14[21]);
FA1A GS14_22(ps15[21], pc15[22], g14[22], ps14[22], pc14[22]);
FA1A GS14_23(ps15[22], pc15[23], g14[23], ps14[23], pc14[23]);
FA1A GS14_24(ps15[23], pc15[24], g14[24], ps14[24], pc14[24]);
FA1A GS14_25(ps15[24], pc15[25], g14[25], ps14[25], pc14[25]);
FA1A GS14_26(ps15[25], pc15[26], g14[26], ps14[26], pc14[26]);
FA1A GS14_27(ps15[26], pc15[27], g14[27], ps14[27], pc14[27]);
FA1A GS14_28(ps15[27], pc15[28], g14[28], ps14[28], pc14[28]);
FA1A GS14_29(ps15[28], pc15[29], g14[29], ps14[29], pc14[29]);
FA1A GS14_30(ps15[29], pc15[30], g14[30], ps14[30], pc14[30]);
FA1A GS14_31(ps15[30], pc15[31], g14[31], ps14[31], pc14[31]);
FA1A GS14_32(ps15[31], pc15[32], g14[32], ps14[32], pc14[32]);
FA1A GS14_33(ps15[32], pc15[33], g14[33], ps14[33], pc14[33]);
FA1A GS14_34(ps15[33], pc15[34], g14[34], ps14[34], pc14[34]);
FA1A GS14_35(ps15[34], pc15[35], g14[35], ps14[35], pc14[35]);
FA1A GS14_36(ps15[35], pc15[36], g14[36], ps14[36], pc14[36]);
FA1A GS14_37(ps15[36], pc15[37], g14[37], ps14[37], pc14[37]);
FA1A GS14_38(ps15[37], pc15[38], g14[38], ps14[38], pc14[38]);
FA1A GS14_39(ps15[38], pc15[39], g14[39], ps14[39], pc14[39]);
FA1A GS14_40(ps15[39], pc15[40], g14[40], ps14[40], pc14[40]);
FA1A GS14_41(ps15[40], pc15[41], g14[41], ps14[41], pc14[41]);
FA1A GS14_42(ps15[41], pc15[42], g14[42], ps14[42], pc14[42]);
FA1A GS14_43(ps15[42], pc15[43], g14[43], ps14[43], pc14[43]);
FA1A GS14_44(ps15[43], pc15[44], g14[44], ps14[44], pc14[44]);
FA1A GS14_45(ps15[44], pc15[45], g14[45], ps14[45], pc14[45]);
FA1A GS14_46(ps15[45], pc15[46], g14[46], ps14[46], pc14[46]);
FA1A GS14_47(ps15[46], pc15[47], g14[47], ps14[47], pc14[47]);
FA1A GS14_48(ps15[47], pc15[48], g14[48], ps14[48], pc14[48]);
FA1A GS14_49(ps15[48], pc15[49], g14[49], ps14[49], pc14[49]);
FA1A GS14_50(ps15[49], pc15[50], g14[50], ps14[50], pc14[50]);
FA1A GS14_51(ps15[50], pc15[51], g14[51], ps14[51], pc14[51]);
FA1A GS14_52(ps15[51], pc15[52], g14[52], ps14[52], pc14[52]);
FA1A GS14_53(ps15[52], pc15[53], g14[53], ps14[53], pc14[53]);
FA1A GS14_54(ps15[53], pc15[54], g14[54], ps14[54], pc14[54]);
FA1A GS14_55(ps15[54], pc15[55], g14[55], ps14[55], pc14[55]);
FA1A GS14_56(ps15[55], pc15[56], g14[56], ps14[56], pc14[56]);
FA1A GS14_57(ps15[56], pc15[57], g14[57], ps14[57], pc14[57]);
FA1A GS14_58(ps15[57], pc15[58], g14[58], ps14[58], pc14[58]);
FA1A GS14_59(ps15[58], pc15[59], g14[59], ps14[59], pc14[59]);
FA1A GS14_60(ps15[59], pc15[60], g14[60], ps14[60], pc14[60]);
FA1A GS14_61(ps15[60], pc15[61], g14[61], ps14[61], pc14[61]);
FA1A GS14_62(ps15[61], pc15[62], g14[62], ps14[62], pc14[62]);
FA1A GS14_63(ps15[62], pc15[63], g14[63], ps14[63], pc14[63]);
FA1A GS13_9(g14[8], pc14[9], g13[9], ps13[9], pc13[9]);
FA1A GS13_10(ps14[9], pc14[10], g13[10], ps13[10], pc13[10]);
FA1A GS13_11(ps14[10], pc14[11], g13[11], ps13[11], pc13[11]);
FA1A GS13_12(ps14[11], pc14[12], g13[12], ps13[12], pc13[12]);
FA1A GS13_13(ps14[12], pc14[13], g13[13], ps13[13], pc13[13]);
FA1A GS13_14(ps14[13], pc14[14], g13[14], ps13[14], pc13[14]);
FA1A GS13_15(ps14[14], pc14[15], g13[15], ps13[15], pc13[15]);
FA1A GS13_16(ps14[15], pc14[16], g13[16], ps13[16], pc13[16]);
FA1A GS13_17(ps14[16], pc14[17], g13[17], ps13[17], pc13[17]);
FA1A GS13_18(ps14[17], pc14[18], g13[18], ps13[18], pc13[18]);
FA1A GS13_19(ps14[18], pc14[19], g13[19], ps13[19], pc13[19]);
FA1A GS13_20(ps14[19], pc14[20], g13[20], ps13[20], pc13[20]);
FA1A GS13_21(ps14[20], pc14[21], g13[21], ps13[21], pc13[21]);
FA1A GS13_22(ps14[21], pc14[22], g13[22], ps13[22], pc13[22]);
FA1A GS13_23(ps14[22], pc14[23], g13[23], ps13[23], pc13[23]);
FA1A GS13_24(ps14[23], pc14[24], g13[24], ps13[24], pc13[24]);
FA1A GS13_25(ps14[24], pc14[25], g13[25], ps13[25], pc13[25]);
FA1A GS13_26(ps14[25], pc14[26], g13[26], ps13[26], pc13[26]);
FA1A GS13_27(ps14[26], pc14[27], g13[27], ps13[27], pc13[27]);
FA1A GS13_28(ps14[27], pc14[28], g13[28], ps13[28], pc13[28]);
FA1A GS13_29(ps14[28], pc14[29], g13[29], ps13[29], pc13[29]);
FA1A GS13_30(ps14[29], pc14[30], g13[30], ps13[30], pc13[30]);
FA1A GS13_31(ps14[30], pc14[31], g13[31], ps13[31], pc13[31]);
FA1A GS13_32(ps14[31], pc14[32], g13[32], ps13[32], pc13[32]);
FA1A GS13_33(ps14[32], pc14[33], g13[33], ps13[33], pc13[33]);
FA1A GS13_34(ps14[33], pc14[34], g13[34], ps13[34], pc13[34]);
FA1A GS13_35(ps14[34], pc14[35], g13[35], ps13[35], pc13[35]);
FA1A GS13_36(ps14[35], pc14[36], g13[36], ps13[36], pc13[36]);
FA1A GS13_37(ps14[36], pc14[37], g13[37], ps13[37], pc13[37]);
FA1A GS13_38(ps14[37], pc14[38], g13[38], ps13[38], pc13[38]);
FA1A GS13_39(ps14[38], pc14[39], g13[39], ps13[39], pc13[39]);
FA1A GS13_40(ps14[39], pc14[40], g13[40], ps13[40], pc13[40]);
FA1A GS13_41(ps14[40], pc14[41], g13[41], ps13[41], pc13[41]);
FA1A GS13_42(ps14[41], pc14[42], g13[42], ps13[42], pc13[42]);
FA1A GS13_43(ps14[42], pc14[43], g13[43], ps13[43], pc13[43]);
FA1A GS13_44(ps14[43], pc14[44], g13[44], ps13[44], pc13[44]);
FA1A GS13_45(ps14[44], pc14[45], g13[45], ps13[45], pc13[45]);
FA1A GS13_46(ps14[45], pc14[46], g13[46], ps13[46], pc13[46]);
FA1A GS13_47(ps14[46], pc14[47], g13[47], ps13[47], pc13[47]);
FA1A GS13_48(ps14[47], pc14[48], g13[48], ps13[48], pc13[48]);
FA1A GS13_49(ps14[48], pc14[49], g13[49], ps13[49], pc13[49]);
FA1A GS13_50(ps14[49], pc14[50], g13[50], ps13[50], pc13[50]);
FA1A GS13_51(ps14[50], pc14[51], g13[51], ps13[51], pc13[51]);
FA1A GS13_52(ps14[51], pc14[52], g13[52], ps13[52], pc13[52]);
FA1A GS13_53(ps14[52], pc14[53], g13[53], ps13[53], pc13[53]);
FA1A GS13_54(ps14[53], pc14[54], g13[54], ps13[54], pc13[54]);
FA1A GS13_55(ps14[54], pc14[55], g13[55], ps13[55], pc13[55]);
FA1A GS13_56(ps14[55], pc14[56], g13[56], ps13[56], pc13[56]);
FA1A GS13_57(ps14[56], pc14[57], g13[57], ps13[57], pc13[57]);
FA1A GS13_58(ps14[57], pc14[58], g13[58], ps13[58], pc13[58]);
FA1A GS13_59(ps14[58], pc14[59], g13[59], ps13[59], pc13[59]);
FA1A GS13_60(ps14[59], pc14[60], g13[60], ps13[60], pc13[60]);
FA1A GS13_61(ps14[60], pc14[61], g13[61], ps13[61], pc13[61]);
FA1A GS13_62(ps14[61], pc14[62], g13[62], ps13[62], pc13[62]);
FA1A GS13_63(ps14[62], pc14[63], g13[63], ps13[63], pc13[63]);
FA1A GS12_9(g13[8], pc13[9], g12[9], ps12[9], pc12[9]);
FA1A GS12_10(ps13[9], pc13[10], g12[10], ps12[10], pc12[10]);
FA1A GS12_11(ps13[10], pc13[11], g12[11], ps12[11], pc12[11]);
FA1A GS12_12(ps13[11], pc13[12], g12[12], ps12[12], pc12[12]);
FA1A GS12_13(ps13[12], pc13[13], g12[13], ps12[13], pc12[13]);
FA1A GS12_14(ps13[13], pc13[14], g12[14], ps12[14], pc12[14]);
FA1A GS12_15(ps13[14], pc13[15], g12[15], ps12[15], pc12[15]);
FA1A GS12_16(ps13[15], pc13[16], g12[16], ps12[16], pc12[16]);
FA1A GS12_17(ps13[16], pc13[17], g12[17], ps12[17], pc12[17]);
FA1A GS12_18(ps13[17], pc13[18], g12[18], ps12[18], pc12[18]);
FA1A GS12_19(ps13[18], pc13[19], g12[19], ps12[19], pc12[19]);
FA1A GS12_20(ps13[19], pc13[20], g12[20], ps12[20], pc12[20]);
FA1A GS12_21(ps13[20], pc13[21], g12[21], ps12[21], pc12[21]);
FA1A GS12_22(ps13[21], pc13[22], g12[22], ps12[22], pc12[22]);
FA1A GS12_23(ps13[22], pc13[23], g12[23], ps12[23], pc12[23]);
FA1A GS12_24(ps13[23], pc13[24], g12[24], ps12[24], pc12[24]);
FA1A GS12_25(ps13[24], pc13[25], g12[25], ps12[25], pc12[25]);
FA1A GS12_26(ps13[25], pc13[26], g12[26], ps12[26], pc12[26]);
FA1A GS12_27(ps13[26], pc13[27], g12[27], ps12[27], pc12[27]);
FA1A GS12_28(ps13[27], pc13[28], g12[28], ps12[28], pc12[28]);
FA1A GS12_29(ps13[28], pc13[29], g12[29], ps12[29], pc12[29]);
FA1A GS12_30(ps13[29], pc13[30], g12[30], ps12[30], pc12[30]);
FA1A GS12_31(ps13[30], pc13[31], g12[31], ps12[31], pc12[31]);
FA1A GS12_32(ps13[31], pc13[32], g12[32], ps12[32], pc12[32]);
FA1A GS12_33(ps13[32], pc13[33], g12[33], ps12[33], pc12[33]);
FA1A GS12_34(ps13[33], pc13[34], g12[34], ps12[34], pc12[34]);
FA1A GS12_35(ps13[34], pc13[35], g12[35], ps12[35], pc12[35]);
FA1A GS12_36(ps13[35], pc13[36], g12[36], ps12[36], pc12[36]);
FA1A GS12_37(ps13[36], pc13[37], g12[37], ps12[37], pc12[37]);
FA1A GS12_38(ps13[37], pc13[38], g12[38], ps12[38], pc12[38]);
FA1A GS12_39(ps13[38], pc13[39], g12[39], ps12[39], pc12[39]);
FA1A GS12_40(ps13[39], pc13[40], g12[40], ps12[40], pc12[40]);
FA1A GS12_41(ps13[40], pc13[41], g12[41], ps12[41], pc12[41]);
FA1A GS12_42(ps13[41], pc13[42], g12[42], ps12[42], pc12[42]);
FA1A GS12_43(ps13[42], pc13[43], g12[43], ps12[43], pc12[43]);
FA1A GS12_44(ps13[43], pc13[44], g12[44], ps12[44], pc12[44]);
FA1A GS12_45(ps13[44], pc13[45], g12[45], ps12[45], pc12[45]);
FA1A GS12_46(ps13[45], pc13[46], g12[46], ps12[46], pc12[46]);
FA1A GS12_47(ps13[46], pc13[47], g12[47], ps12[47], pc12[47]);
FA1A GS12_48(ps13[47], pc13[48], g12[48], ps12[48], pc12[48]);
FA1A GS12_49(ps13[48], pc13[49], g12[49], ps12[49], pc12[49]);
FA1A GS12_50(ps13[49], pc13[50], g12[50], ps12[50], pc12[50]);
FA1A GS12_51(ps13[50], pc13[51], g12[51], ps12[51], pc12[51]);
FA1A GS12_52(ps13[51], pc13[52], g12[52], ps12[52], pc12[52]);
FA1A GS12_53(ps13[52], pc13[53], g12[53], ps12[53], pc12[53]);
FA1A GS12_54(ps13[53], pc13[54], g12[54], ps12[54], pc12[54]);
FA1A GS12_55(ps13[54], pc13[55], g12[55], ps12[55], pc12[55]);
FA1A GS12_56(ps13[55], pc13[56], g12[56], ps12[56], pc12[56]);
FA1A GS12_57(ps13[56], pc13[57], g12[57], ps12[57], pc12[57]);
FA1A GS12_58(ps13[57], pc13[58], g12[58], ps12[58], pc12[58]);
FA1A GS12_59(ps13[58], pc13[59], g12[59], ps12[59], pc12[59]);
FA1A GS12_60(ps13[59], pc13[60], g12[60], ps12[60], pc12[60]);
FA1A GS12_61(ps13[60], pc13[61], g12[61], ps12[61], pc12[61]);
FA1A GS12_62(ps13[61], pc13[62], g12[62], ps12[62], pc12[62]);
FA1A GS12_63(ps13[62], pc13[63], g12[63], ps12[63], pc12[63]);
FA1A GS11_9(g12[8], pc12[9], g11[9], ps11[9], pc11[9]);
FA1A GS11_10(ps12[9], pc12[10], g11[10], ps11[10], pc11[10]);
FA1A GS11_11(ps12[10], pc12[11], g11[11], ps11[11], pc11[11]);
FA1A GS11_12(ps12[11], pc12[12], g11[12], ps11[12], pc11[12]);
FA1A GS11_13(ps12[12], pc12[13], g11[13], ps11[13], pc11[13]);
FA1A GS11_14(ps12[13], pc12[14], g11[14], ps11[14], pc11[14]);
FA1A GS11_15(ps12[14], pc12[15], g11[15], ps11[15], pc11[15]);
FA1A GS11_16(ps12[15], pc12[16], g11[16], ps11[16], pc11[16]);
FA1A GS11_17(ps12[16], pc12[17], g11[17], ps11[17], pc11[17]);
FA1A GS11_18(ps12[17], pc12[18], g11[18], ps11[18], pc11[18]);
FA1A GS11_19(ps12[18], pc12[19], g11[19], ps11[19], pc11[19]);
FA1A GS11_20(ps12[19], pc12[20], g11[20], ps11[20], pc11[20]);
FA1A GS11_21(ps12[20], pc12[21], g11[21], ps11[21], pc11[21]);
FA1A GS11_22(ps12[21], pc12[22], g11[22], ps11[22], pc11[22]);
FA1A GS11_23(ps12[22], pc12[23], g11[23], ps11[23], pc11[23]);
FA1A GS11_24(ps12[23], pc12[24], g11[24], ps11[24], pc11[24]);
FA1A GS11_25(ps12[24], pc12[25], g11[25], ps11[25], pc11[25]);
FA1A GS11_26(ps12[25], pc12[26], g11[26], ps11[26], pc11[26]);
FA1A GS11_27(ps12[26], pc12[27], g11[27], ps11[27], pc11[27]);
FA1A GS11_28(ps12[27], pc12[28], g11[28], ps11[28], pc11[28]);
FA1A GS11_29(ps12[28], pc12[29], g11[29], ps11[29], pc11[29]);
FA1A GS11_30(ps12[29], pc12[30], g11[30], ps11[30], pc11[30]);
FA1A GS11_31(ps12[30], pc12[31], g11[31], ps11[31], pc11[31]);
FA1A GS11_32(ps12[31], pc12[32], g11[32], ps11[32], pc11[32]);
FA1A GS11_33(ps12[32], pc12[33], g11[33], ps11[33], pc11[33]);
FA1A GS11_34(ps12[33], pc12[34], g11[34], ps11[34], pc11[34]);
FA1A GS11_35(ps12[34], pc12[35], g11[35], ps11[35], pc11[35]);
FA1A GS11_36(ps12[35], pc12[36], g11[36], ps11[36], pc11[36]);
FA1A GS11_37(ps12[36], pc12[37], g11[37], ps11[37], pc11[37]);
FA1A GS11_38(ps12[37], pc12[38], g11[38], ps11[38], pc11[38]);
FA1A GS11_39(ps12[38], pc12[39], g11[39], ps11[39], pc11[39]);
FA1A GS11_40(ps12[39], pc12[40], g11[40], ps11[40], pc11[40]);
FA1A GS11_41(ps12[40], pc12[41], g11[41], ps11[41], pc11[41]);
FA1A GS11_42(ps12[41], pc12[42], g11[42], ps11[42], pc11[42]);
FA1A GS11_43(ps12[42], pc12[43], g11[43], ps11[43], pc11[43]);
FA1A GS11_44(ps12[43], pc12[44], g11[44], ps11[44], pc11[44]);
FA1A GS11_45(ps12[44], pc12[45], g11[45], ps11[45], pc11[45]);
FA1A GS11_46(ps12[45], pc12[46], g11[46], ps11[46], pc11[46]);
FA1A GS11_47(ps12[46], pc12[47], g11[47], ps11[47], pc11[47]);
FA1A GS11_48(ps12[47], pc12[48], g11[48], ps11[48], pc11[48]);
FA1A GS11_49(ps12[48], pc12[49], g11[49], ps11[49], pc11[49]);
FA1A GS11_50(ps12[49], pc12[50], g11[50], ps11[50], pc11[50]);
FA1A GS11_51(ps12[50], pc12[51], g11[51], ps11[51], pc11[51]);
FA1A GS11_52(ps12[51], pc12[52], g11[52], ps11[52], pc11[52]);
FA1A GS11_53(ps12[52], pc12[53], g11[53], ps11[53], pc11[53]);
FA1A GS11_54(ps12[53], pc12[54], g11[54], ps11[54], pc11[54]);
FA1A GS11_55(ps12[54], pc12[55], g11[55], ps11[55], pc11[55]);
FA1A GS11_56(ps12[55], pc12[56], g11[56], ps11[56], pc11[56]);
FA1A GS11_57(ps12[56], pc12[57], g11[57], ps11[57], pc11[57]);
FA1A GS11_58(ps12[57], pc12[58], g11[58], ps11[58], pc11[58]);
FA1A GS11_59(ps12[58], pc12[59], g11[59], ps11[59], pc11[59]);
FA1A GS11_60(ps12[59], pc12[60], g11[60], ps11[60], pc11[60]);
FA1A GS11_61(ps12[60], pc12[61], g11[61], ps11[61], pc11[61]);
FA1A GS11_62(ps12[61], pc12[62], g11[62], ps11[62], pc11[62]);
FA1A GS11_63(ps12[62], pc12[63], g11[63], ps11[63], pc11[63]);
FA1A GS10_9(g11[8], pc11[9], g10[9], ps10[9], pc10[9]);
FA1A GS10_10(ps11[9], pc11[10], g10[10], ps10[10], pc10[10]);
FA1A GS10_11(ps11[10], pc11[11], g10[11], ps10[11], pc10[11]);
FA1A GS10_12(ps11[11], pc11[12], g10[12], ps10[12], pc10[12]);
FA1A GS10_13(ps11[12], pc11[13], g10[13], ps10[13], pc10[13]);
FA1A GS10_14(ps11[13], pc11[14], g10[14], ps10[14], pc10[14]);
FA1A GS10_15(ps11[14], pc11[15], g10[15], ps10[15], pc10[15]);
FA1A GS10_16(ps11[15], pc11[16], g10[16], ps10[16], pc10[16]);
FA1A GS10_17(ps11[16], pc11[17], g10[17], ps10[17], pc10[17]);
FA1A GS10_18(ps11[17], pc11[18], g10[18], ps10[18], pc10[18]);
FA1A GS10_19(ps11[18], pc11[19], g10[19], ps10[19], pc10[19]);
FA1A GS10_20(ps11[19], pc11[20], g10[20], ps10[20], pc10[20]);
FA1A GS10_21(ps11[20], pc11[21], g10[21], ps10[21], pc10[21]);
FA1A GS10_22(ps11[21], pc11[22], g10[22], ps10[22], pc10[22]);
FA1A GS10_23(ps11[22], pc11[23], g10[23], ps10[23], pc10[23]);
FA1A GS10_24(ps11[23], pc11[24], g10[24], ps10[24], pc10[24]);
FA1A GS10_25(ps11[24], pc11[25], g10[25], ps10[25], pc10[25]);
FA1A GS10_26(ps11[25], pc11[26], g10[26], ps10[26], pc10[26]);
FA1A GS10_27(ps11[26], pc11[27], g10[27], ps10[27], pc10[27]);
FA1A GS10_28(ps11[27], pc11[28], g10[28], ps10[28], pc10[28]);
FA1A GS10_29(ps11[28], pc11[29], g10[29], ps10[29], pc10[29]);
FA1A GS10_30(ps11[29], pc11[30], g10[30], ps10[30], pc10[30]);
FA1A GS10_31(ps11[30], pc11[31], g10[31], ps10[31], pc10[31]);
FA1A GS10_32(ps11[31], pc11[32], g10[32], ps10[32], pc10[32]);
FA1A GS10_33(ps11[32], pc11[33], g10[33], ps10[33], pc10[33]);
FA1A GS10_34(ps11[33], pc11[34], g10[34], ps10[34], pc10[34]);
FA1A GS10_35(ps11[34], pc11[35], g10[35], ps10[35], pc10[35]);
FA1A GS10_36(ps11[35], pc11[36], g10[36], ps10[36], pc10[36]);
FA1A GS10_37(ps11[36], pc11[37], g10[37], ps10[37], pc10[37]);
FA1A GS10_38(ps11[37], pc11[38], g10[38], ps10[38], pc10[38]);
FA1A GS10_39(ps11[38], pc11[39], g10[39], ps10[39], pc10[39]);
FA1A GS10_40(ps11[39], pc11[40], g10[40], ps10[40], pc10[40]);
FA1A GS10_41(ps11[40], pc11[41], g10[41], ps10[41], pc10[41]);
FA1A GS10_42(ps11[41], pc11[42], g10[42], ps10[42], pc10[42]);
FA1A GS10_43(ps11[42], pc11[43], g10[43], ps10[43], pc10[43]);
FA1A GS10_44(ps11[43], pc11[44], g10[44], ps10[44], pc10[44]);
FA1A GS10_45(ps11[44], pc11[45], g10[45], ps10[45], pc10[45]);
FA1A GS10_46(ps11[45], pc11[46], g10[46], ps10[46], pc10[46]);
FA1A GS10_47(ps11[46], pc11[47], g10[47], ps10[47], pc10[47]);
FA1A GS10_48(ps11[47], pc11[48], g10[48], ps10[48], pc10[48]);
FA1A GS10_49(ps11[48], pc11[49], g10[49], ps10[49], pc10[49]);
FA1A GS10_50(ps11[49], pc11[50], g10[50], ps10[50], pc10[50]);
FA1A GS10_51(ps11[50], pc11[51], g10[51], ps10[51], pc10[51]);
FA1A GS10_52(ps11[51], pc11[52], g10[52], ps10[52], pc10[52]);
FA1A GS10_53(ps11[52], pc11[53], g10[53], ps10[53], pc10[53]);
FA1A GS10_54(ps11[53], pc11[54], g10[54], ps10[54], pc10[54]);
FA1A GS10_55(ps11[54], pc11[55], g10[55], ps10[55], pc10[55]);
FA1A GS10_56(ps11[55], pc11[56], g10[56], ps10[56], pc10[56]);
FA1A GS10_57(ps11[56], pc11[57], g10[57], ps10[57], pc10[57]);
FA1A GS10_58(ps11[57], pc11[58], g10[58], ps10[58], pc10[58]);
FA1A GS10_59(ps11[58], pc11[59], g10[59], ps10[59], pc10[59]);
FA1A GS10_60(ps11[59], pc11[60], g10[60], ps10[60], pc10[60]);
FA1A GS10_61(ps11[60], pc11[61], g10[61], ps10[61], pc10[61]);
FA1A GS10_62(ps11[61], pc11[62], g10[62], ps10[62], pc10[62]);
FA1A GS10_63(ps11[62], pc11[63], g10[63], ps10[63], pc10[63]);
FA1A GS9_9(g10[8], pc10[9], g9[9], ps9[9], pc9[9]);
FA1A GS9_10(ps10[9], pc10[10], g9[10], ps9[10], pc9[10]);
FA1A GS9_11(ps10[10], pc10[11], g9[11], ps9[11], pc9[11]);
FA1A GS9_12(ps10[11], pc10[12], g9[12], ps9[12], pc9[12]);
FA1A GS9_13(ps10[12], pc10[13], g9[13], ps9[13], pc9[13]);
FA1A GS9_14(ps10[13], pc10[14], g9[14], ps9[14], pc9[14]);
FA1A GS9_15(ps10[14], pc10[15], g9[15], ps9[15], pc9[15]);
FA1A GS9_16(ps10[15], pc10[16], g9[16], ps9[16], pc9[16]);
FA1A GS9_17(ps10[16], pc10[17], g9[17], ps9[17], pc9[17]);
FA1A GS9_18(ps10[17], pc10[18], g9[18], ps9[18], pc9[18]);
FA1A GS9_19(ps10[18], pc10[19], g9[19], ps9[19], pc9[19]);
FA1A GS9_20(ps10[19], pc10[20], g9[20], ps9[20], pc9[20]);
FA1A GS9_21(ps10[20], pc10[21], g9[21], ps9[21], pc9[21]);
FA1A GS9_22(ps10[21], pc10[22], g9[22], ps9[22], pc9[22]);
FA1A GS9_23(ps10[22], pc10[23], g9[23], ps9[23], pc9[23]);
FA1A GS9_24(ps10[23], pc10[24], g9[24], ps9[24], pc9[24]);
FA1A GS9_25(ps10[24], pc10[25], g9[25], ps9[25], pc9[25]);
FA1A GS9_26(ps10[25], pc10[26], g9[26], ps9[26], pc9[26]);
FA1A GS9_27(ps10[26], pc10[27], g9[27], ps9[27], pc9[27]);
FA1A GS9_28(ps10[27], pc10[28], g9[28], ps9[28], pc9[28]);
FA1A GS9_29(ps10[28], pc10[29], g9[29], ps9[29], pc9[29]);
FA1A GS9_30(ps10[29], pc10[30], g9[30], ps9[30], pc9[30]);
FA1A GS9_31(ps10[30], pc10[31], g9[31], ps9[31], pc9[31]);
FA1A GS9_32(ps10[31], pc10[32], g9[32], ps9[32], pc9[32]);
FA1A GS9_33(ps10[32], pc10[33], g9[33], ps9[33], pc9[33]);
FA1A GS9_34(ps10[33], pc10[34], g9[34], ps9[34], pc9[34]);
FA1A GS9_35(ps10[34], pc10[35], g9[35], ps9[35], pc9[35]);
FA1A GS9_36(ps10[35], pc10[36], g9[36], ps9[36], pc9[36]);
FA1A GS9_37(ps10[36], pc10[37], g9[37], ps9[37], pc9[37]);
FA1A GS9_38(ps10[37], pc10[38], g9[38], ps9[38], pc9[38]);
FA1A GS9_39(ps10[38], pc10[39], g9[39], ps9[39], pc9[39]);
FA1A GS9_40(ps10[39], pc10[40], g9[40], ps9[40], pc9[40]);
FA1A GS9_41(ps10[40], pc10[41], g9[41], ps9[41], pc9[41]);
FA1A GS9_42(ps10[41], pc10[42], g9[42], ps9[42], pc9[42]);
FA1A GS9_43(ps10[42], pc10[43], g9[43], ps9[43], pc9[43]);
FA1A GS9_44(ps10[43], pc10[44], g9[44], ps9[44], pc9[44]);
FA1A GS9_45(ps10[44], pc10[45], g9[45], ps9[45], pc9[45]);
FA1A GS9_46(ps10[45], pc10[46], g9[46], ps9[46], pc9[46]);
FA1A GS9_47(ps10[46], pc10[47], g9[47], ps9[47], pc9[47]);
FA1A GS9_48(ps10[47], pc10[48], g9[48], ps9[48], pc9[48]);
FA1A GS9_49(ps10[48], pc10[49], g9[49], ps9[49], pc9[49]);
FA1A GS9_50(ps10[49], pc10[50], g9[50], ps9[50], pc9[50]);
FA1A GS9_51(ps10[50], pc10[51], g9[51], ps9[51], pc9[51]);
FA1A GS9_52(ps10[51], pc10[52], g9[52], ps9[52], pc9[52]);
FA1A GS9_53(ps10[52], pc10[53], g9[53], ps9[53], pc9[53]);
FA1A GS9_54(ps10[53], pc10[54], g9[54], ps9[54], pc9[54]);
FA1A GS9_55(ps10[54], pc10[55], g9[55], ps9[55], pc9[55]);
FA1A GS9_56(ps10[55], pc10[56], g9[56], ps9[56], pc9[56]);
FA1A GS9_57(ps10[56], pc10[57], g9[57], ps9[57], pc9[57]);
FA1A GS9_58(ps10[57], pc10[58], g9[58], ps9[58], pc9[58]);
FA1A GS9_59(ps10[58], pc10[59], g9[59], ps9[59], pc9[59]);
FA1A GS9_60(ps10[59], pc10[60], g9[60], ps9[60], pc9[60]);
FA1A GS9_61(ps10[60], pc10[61], g9[61], ps9[61], pc9[61]);
FA1A GS9_62(ps10[61], pc10[62], g9[62], ps9[62], pc9[62]);
FA1A GS9_63(ps10[62], pc10[63], g9[63], ps9[63], pc9[63]);
FA1A GS8_9(g9[8], pc9[9], g8[9], ps8[9], pc8[9]);
FA1A GS8_10(ps9[9], pc9[10], g8[10], ps8[10], pc8[10]);
FA1A GS8_11(ps9[10], pc9[11], g8[11], ps8[11], pc8[11]);
FA1A GS8_12(ps9[11], pc9[12], g8[12], ps8[12], pc8[12]);
FA1A GS8_13(ps9[12], pc9[13], g8[13], ps8[13], pc8[13]);
FA1A GS8_14(ps9[13], pc9[14], g8[14], ps8[14], pc8[14]);
FA1A GS8_15(ps9[14], pc9[15], g8[15], ps8[15], pc8[15]);
FA1A GS8_16(ps9[15], pc9[16], g8[16], ps8[16], pc8[16]);
FA1A GS8_17(ps9[16], pc9[17], g8[17], ps8[17], pc8[17]);
FA1A GS8_18(ps9[17], pc9[18], g8[18], ps8[18], pc8[18]);
FA1A GS8_19(ps9[18], pc9[19], g8[19], ps8[19], pc8[19]);
FA1A GS8_20(ps9[19], pc9[20], g8[20], ps8[20], pc8[20]);
FA1A GS8_21(ps9[20], pc9[21], g8[21], ps8[21], pc8[21]);
FA1A GS8_22(ps9[21], pc9[22], g8[22], ps8[22], pc8[22]);
FA1A GS8_23(ps9[22], pc9[23], g8[23], ps8[23], pc8[23]);
FA1A GS8_24(ps9[23], pc9[24], g8[24], ps8[24], pc8[24]);
FA1A GS8_25(ps9[24], pc9[25], g8[25], ps8[25], pc8[25]);
FA1A GS8_26(ps9[25], pc9[26], g8[26], ps8[26], pc8[26]);
FA1A GS8_27(ps9[26], pc9[27], g8[27], ps8[27], pc8[27]);
FA1A GS8_28(ps9[27], pc9[28], g8[28], ps8[28], pc8[28]);
FA1A GS8_29(ps9[28], pc9[29], g8[29], ps8[29], pc8[29]);
FA1A GS8_30(ps9[29], pc9[30], g8[30], ps8[30], pc8[30]);
FA1A GS8_31(ps9[30], pc9[31], g8[31], ps8[31], pc8[31]);
FA1A GS8_32(ps9[31], pc9[32], g8[32], ps8[32], pc8[32]);
FA1A GS8_33(ps9[32], pc9[33], g8[33], ps8[33], pc8[33]);
FA1A GS8_34(ps9[33], pc9[34], g8[34], ps8[34], pc8[34]);
FA1A GS8_35(ps9[34], pc9[35], g8[35], ps8[35], pc8[35]);
FA1A GS8_36(ps9[35], pc9[36], g8[36], ps8[36], pc8[36]);
FA1A GS8_37(ps9[36], pc9[37], g8[37], ps8[37], pc8[37]);
FA1A GS8_38(ps9[37], pc9[38], g8[38], ps8[38], pc8[38]);
FA1A GS8_39(ps9[38], pc9[39], g8[39], ps8[39], pc8[39]);
FA1A GS8_40(ps9[39], pc9[40], g8[40], ps8[40], pc8[40]);
FA1A GS8_41(ps9[40], pc9[41], g8[41], ps8[41], pc8[41]);
FA1A GS8_42(ps9[41], pc9[42], g8[42], ps8[42], pc8[42]);
FA1A GS8_43(ps9[42], pc9[43], g8[43], ps8[43], pc8[43]);
FA1A GS8_44(ps9[43], pc9[44], g8[44], ps8[44], pc8[44]);
FA1A GS8_45(ps9[44], pc9[45], g8[45], ps8[45], pc8[45]);
FA1A GS8_46(ps9[45], pc9[46], g8[46], ps8[46], pc8[46]);
FA1A GS8_47(ps9[46], pc9[47], g8[47], ps8[47], pc8[47]);
FA1A GS8_48(ps9[47], pc9[48], g8[48], ps8[48], pc8[48]);
FA1A GS8_49(ps9[48], pc9[49], g8[49], ps8[49], pc8[49]);
FA1A GS8_50(ps9[49], pc9[50], g8[50], ps8[50], pc8[50]);
FA1A GS8_51(ps9[50], pc9[51], g8[51], ps8[51], pc8[51]);
FA1A GS8_52(ps9[51], pc9[52], g8[52], ps8[52], pc8[52]);
FA1A GS8_53(ps9[52], pc9[53], g8[53], ps8[53], pc8[53]);
FA1A GS8_54(ps9[53], pc9[54], g8[54], ps8[54], pc8[54]);
FA1A GS8_55(ps9[54], pc9[55], g8[55], ps8[55], pc8[55]);
FA1A GS8_56(ps9[55], pc9[56], g8[56], ps8[56], pc8[56]);
FA1A GS8_57(ps9[56], pc9[57], g8[57], ps8[57], pc8[57]);
FA1A GS8_58(ps9[57], pc9[58], g8[58], ps8[58], pc8[58]);
FA1A GS8_59(ps9[58], pc9[59], g8[59], ps8[59], pc8[59]);
FA1A GS8_60(ps9[59], pc9[60], g8[60], ps8[60], pc8[60]);
FA1A GS8_61(ps9[60], pc9[61], g8[61], ps8[61], pc8[61]);
FA1A GS8_62(ps9[61], pc9[62], g8[62], ps8[62], pc8[62]);
FA1A GS8_63(ps9[62], pc9[63], g8[63], product[63], pc8[63]);
AN2 GANDG_8(g8[8], pc8[9], gen[8]);
AN2 GANDG_9(ps8[9], pc8[10], gen[9]);
AN2 GANDG_10(ps8[10], pc8[11], gen[10]);
AN2 GANDG_11(ps8[11], pc8[12], gen[11]);
AN2 GANDG_12(ps8[12], pc8[13], gen[12]);
AN2 GANDG_13(ps8[13], pc8[14], gen[13]);
AN2 GANDG_14(ps8[14], pc8[15], gen[14]);
AN2 GANDG_15(ps8[15], pc8[16], gen[15]);
AN2 GANDG_16(ps8[16], pc8[17], gen[16]);
AN2 GANDG_17(ps8[17], pc8[18], gen[17]);
AN2 GANDG_18(ps8[18], pc8[19], gen[18]);
AN2 GANDG_19(ps8[19], pc8[20], gen[19]);
AN2 GANDG_20(ps8[20], pc8[21], gen[20]);
AN2 GANDG_21(ps8[21], pc8[22], gen[21]);
AN2 GANDG_22(ps8[22], pc8[23], gen[22]);
AN2 GANDG_23(ps8[23], pc8[24], gen[23]);
AN2 GANDG_24(ps8[24], pc8[25], gen[24]);
AN2 GANDG_25(ps8[25], pc8[26], gen[25]);
AN2 GANDG_26(ps8[26], pc8[27], gen[26]);
AN2 GANDG_27(ps8[27], pc8[28], gen[27]);
AN2 GANDG_28(ps8[28], pc8[29], gen[28]);
AN2 GANDG_29(ps8[29], pc8[30], gen[29]);
AN2 GANDG_30(ps8[30], pc8[31], gen[30]);
AN2 GANDG_31(ps8[31], pc8[32], gen[31]);
AN2 GANDG_32(ps8[32], pc8[33], gen[32]);
AN2 GANDG_33(ps8[33], pc8[34], gen[33]);
AN2 GANDG_34(ps8[34], pc8[35], gen[34]);
AN2 GANDG_35(ps8[35], pc8[36], gen[35]);
AN2 GANDG_36(ps8[36], pc8[37], gen[36]);
AN2 GANDG_37(ps8[37], pc8[38], gen[37]);
AN2 GANDG_38(ps8[38], pc8[39], gen[38]);
AN2 GANDG_39(ps8[39], pc8[40], gen[39]);
AN2 GANDG_40(ps8[40], pc8[41], gen[40]);
AN2 GANDG_41(ps8[41], pc8[42], gen[41]);
AN2 GANDG_42(ps8[42], pc8[43], gen[42]);
AN2 GANDG_43(ps8[43], pc8[44], gen[43]);
AN2 GANDG_44(ps8[44], pc8[45], gen[44]);
AN2 GANDG_45(ps8[45], pc8[46], gen[45]);
AN2 GANDG_46(ps8[46], pc8[47], gen[46]);
AN2 GANDG_47(ps8[47], pc8[48], gen[47]);
AN2 GANDG_48(ps8[48], pc8[49], gen[48]);
AN2 GANDG_49(ps8[49], pc8[50], gen[49]);
AN2 GANDG_50(ps8[50], pc8[51], gen[50]);
AN2 GANDG_51(ps8[51], pc8[52], gen[51]);
AN2 GANDG_52(ps8[52], pc8[53], gen[52]);
AN2 GANDG_53(ps8[53], pc8[54], gen[53]);
AN2 GANDG_54(ps8[54], pc8[55], gen[54]);
AN2 GANDG_55(ps8[55], pc8[56], gen[55]);
AN2 GANDG_56(ps8[56], pc8[57], gen[56]);
AN2 GANDG_57(ps8[57], pc8[58], gen[57]);
AN2 GANDG_58(ps8[58], pc8[59], gen[58]);
AN2 GANDG_59(ps8[59], pc8[60], gen[59]);
AN2 GANDG_60(ps8[60], pc8[61], gen[60]);
AN2 GANDG_61(ps8[61], pc8[62], gen[61]);
AN2 GANDG_62(ps8[62], pc8[63], gen[62]);
OR2 GOR_8(g8[8], pc8[9], tr[8]);
OR2 GOR_9(ps8[9], pc8[10], tr[9]);
OR2 GOR_10(ps8[10], pc8[11], tr[10]);
OR2 GOR_11(ps8[11], pc8[12], tr[11]);
OR2 GOR_12(ps8[12], pc8[13], tr[12]);
OR2 GOR_13(ps8[13], pc8[14], tr[13]);
OR2 GOR_14(ps8[14], pc8[15], tr[14]);
OR2 GOR_15(ps8[15], pc8[16], tr[15]);
OR2 GOR_16(ps8[16], pc8[17], tr[16]);
OR2 GOR_17(ps8[17], pc8[18], tr[17]);
OR2 GOR_18(ps8[18], pc8[19], tr[18]);
OR2 GOR_19(ps8[19], pc8[20], tr[19]);
OR2 GOR_20(ps8[20], pc8[21], tr[20]);
OR2 GOR_21(ps8[21], pc8[22], tr[21]);
OR2 GOR_22(ps8[22], pc8[23], tr[22]);
OR2 GOR_23(ps8[23], pc8[24], tr[23]);
OR2 GOR_24(ps8[24], pc8[25], tr[24]);
OR2 GOR_25(ps8[25], pc8[26], tr[25]);
OR2 GOR_26(ps8[26], pc8[27], tr[26]);
OR2 GOR_27(ps8[27], pc8[28], tr[27]);
OR2 GOR_28(ps8[28], pc8[29], tr[28]);
OR2 GOR_29(ps8[29], pc8[30], tr[29]);
OR2 GOR_30(ps8[30], pc8[31], tr[30]);
OR2 GOR_31(ps8[31], pc8[32], tr[31]);
OR2 GOR_32(ps8[32], pc8[33], tr[32]);
OR2 GOR_33(ps8[33], pc8[34], tr[33]);
OR2 GOR_34(ps8[34], pc8[35], tr[34]);
OR2 GOR_35(ps8[35], pc8[36], tr[35]);
OR2 GOR_36(ps8[36], pc8[37], tr[36]);
OR2 GOR_37(ps8[37], pc8[38], tr[37]);
OR2 GOR_38(ps8[38], pc8[39], tr[38]);
OR2 GOR_39(ps8[39], pc8[40], tr[39]);
OR2 GOR_40(ps8[40], pc8[41], tr[40]);
OR2 GOR_41(ps8[41], pc8[42], tr[41]);
OR2 GOR_42(ps8[42], pc8[43], tr[42]);
OR2 GOR_43(ps8[43], pc8[44], tr[43]);
OR2 GOR_44(ps8[44], pc8[45], tr[44]);
OR2 GOR_45(ps8[45], pc8[46], tr[45]);
OR2 GOR_46(ps8[46], pc8[47], tr[46]);
OR2 GOR_47(ps8[47], pc8[48], tr[47]);
OR2 GOR_48(ps8[48], pc8[49], tr[48]);
OR2 GOR_49(ps8[49], pc8[50], tr[49]);
OR2 GOR_50(ps8[50], pc8[51], tr[50]);
OR2 GOR_51(ps8[51], pc8[52], tr[51]);
OR2 GOR_52(ps8[52], pc8[53], tr[52]);
OR2 GOR_53(ps8[53], pc8[54], tr[53]);
OR2 GOR_54(ps8[54], pc8[55], tr[54]);
OR2 GOR_55(ps8[55], pc8[56], tr[55]);
OR2 GOR_56(ps8[56], pc8[57], tr[56]);
OR2 GOR_57(ps8[57], pc8[58], tr[57]);
OR2 GOR_58(ps8[58], pc8[59], tr[58]);
OR2 GOR_59(ps8[59], pc8[60], tr[59]);
OR2 GOR_60(ps8[60], pc8[61], tr[60]);
OR2 GOR_61(ps8[61], pc8[62], tr[61]);
OR2 GOR_62(ps8[62], pc8[63], tr[62]);
FA1A GFS_8(g8[8], pc8[9], carry[8], product[8], nop[8]);
FA1A GFS_9(ps8[9], pc8[10], carry[9], product[9], nop[9]);
FA1A GFS_10(ps8[10], pc8[11], carry[10], product[10], nop[10]);
FA1A GFS_11(ps8[11], pc8[12], carry[11], product[11], nop[11]);
FA1A GFS_12(ps8[12], pc8[13], carry[12], product[12], nop[12]);
FA1A GFS_13(ps8[13], pc8[14], carry[13], product[13], nop[13]);
FA1A GFS_14(ps8[14], pc8[15], carry[14], product[14], nop[14]);
FA1A GFS_15(ps8[15], pc8[16], carry[15], product[15], nop[15]);
FA1A GFS_16(ps8[16], pc8[17], carry[16], product[16], nop[16]);
FA1A GFS_17(ps8[17], pc8[18], carry[17], product[17], nop[17]);
FA1A GFS_18(ps8[18], pc8[19], carry[18], product[18], nop[18]);
FA1A GFS_19(ps8[19], pc8[20], carry[19], product[19], nop[19]);
FA1A GFS_20(ps8[20], pc8[21], carry[20], product[20], nop[20]);
FA1A GFS_21(ps8[21], pc8[22], carry[21], product[21], nop[21]);
FA1A GFS_22(ps8[22], pc8[23], carry[22], product[22], nop[22]);
FA1A GFS_23(ps8[23], pc8[24], carry[23], product[23], nop[23]);
FA1A GFS_24(ps8[24], pc8[25], carry[24], product[24], nop[24]);
FA1A GFS_25(ps8[25], pc8[26], carry[25], product[25], nop[25]);
FA1A GFS_26(ps8[26], pc8[27], carry[26], product[26], nop[26]);
FA1A GFS_27(ps8[27], pc8[28], carry[27], product[27], nop[27]);
FA1A GFS_28(ps8[28], pc8[29], carry[28], product[28], nop[28]);
FA1A GFS_29(ps8[29], pc8[30], carry[29], product[29], nop[29]);
FA1A GFS_30(ps8[30], pc8[31], carry[30], product[30], nop[30]);
FA1A GFS_31(ps8[31], pc8[32], carry[31], product[31], nop[31]);
FA1A GFS_32(ps8[32], pc8[33], carry[32], product[32], nop[32]);
FA1A GFS_33(ps8[33], pc8[34], carry[33], product[33], nop[33]);
FA1A GFS_34(ps8[34], pc8[35], carry[34], product[34], nop[34]);
FA1A GFS_35(ps8[35], pc8[36], carry[35], product[35], nop[35]);
FA1A GFS_36(ps8[36], pc8[37], carry[36], product[36], nop[36]);
FA1A GFS_37(ps8[37], pc8[38], carry[37], product[37], nop[37]);
FA1A GFS_38(ps8[38], pc8[39], carry[38], product[38], nop[38]);
FA1A GFS_39(ps8[39], pc8[40], carry[39], product[39], nop[39]);
FA1A GFS_40(ps8[40], pc8[41], carry[40], product[40], nop[40]);
FA1A GFS_41(ps8[41], pc8[42], carry[41], product[41], nop[41]);
FA1A GFS_42(ps8[42], pc8[43], carry[42], product[42], nop[42]);
FA1A GFS_43(ps8[43], pc8[44], carry[43], product[43], nop[43]);
FA1A GFS_44(ps8[44], pc8[45], carry[44], product[44], nop[44]);
FA1A GFS_45(ps8[45], pc8[46], carry[45], product[45], nop[45]);
FA1A GFS_46(ps8[46], pc8[47], carry[46], product[46], nop[46]);
FA1A GFS_47(ps8[47], pc8[48], carry[47], product[47], nop[47]);
FA1A GFS_48(ps8[48], pc8[49], carry[48], product[48], nop[48]);
FA1A GFS_49(ps8[49], pc8[50], carry[49], product[49], nop[49]);
FA1A GFS_50(ps8[50], pc8[51], carry[50], product[50], nop[50]);
FA1A GFS_51(ps8[51], pc8[52], carry[51], product[51], nop[51]);
FA1A GFS_52(ps8[52], pc8[53], carry[52], product[52], nop[52]);
FA1A GFS_53(ps8[53], pc8[54], carry[53], product[53], nop[53]);
FA1A GFS_54(ps8[54], pc8[55], carry[54], product[54], nop[54]);
FA1A GFS_55(ps8[55], pc8[56], carry[55], product[55], nop[55]);
FA1A GFS_56(ps8[56], pc8[57], carry[56], product[56], nop[56]);
FA1A GFS_57(ps8[57], pc8[58], carry[57], product[57], nop[57]);
FA1A GFS_58(ps8[58], pc8[59], carry[58], product[58], nop[58]);
FA1A GFS_59(ps8[59], pc8[60], carry[59], product[59], nop[59]);
FA1A GFS_60(ps8[60], pc8[61], carry[60], product[60], nop[60]);
FA1A GFS_61(ps8[61], pc8[62], carry[61], product[61], nop[61]);
FA1A GFS_62(ps8[62], pc8[63], carry[62], product[62], nop[62]);

endmodule

// End of DAS Multiplier circuit


// DA Solutions Ltd., DA Solutions Multiplier/carry block gate level circuit
// Creeated 1-Sep-94, D. J. Wharton
// Circuit also available in VHDL 
// Library used LCA100k CMOS

module carry_block (gen, tr, carry, carry_in, ggen, gtran);

input 	[0:7]	gen, tr;
output 	[0:7]	carry;
input		carry_in;
output		ggen, gtran;

BUF8A CY7(carry_in, carry[7]);
OR2 CY6(gen[7], t76, carry[6]);
AN2 A6A(carry_in, tr[7], t76);
OR3 CY5(gen[6], t75, t65, carry[5]);
AN3 A5A(carry_in, tr[7], tr[6], t75);
AN2 A5B(gen[7], tr[6], t65);
OR4 CY4(gen[5], t74, t64, t54, carry[4]);
AN4 A4A(carry_in, tr[7], tr[6], tr[5], t74);
AN3 A4B(gen[7], tr[6], tr[5], t64);
AN2 A4C(gen[6], tr[5], t54);
OR5 CY3(gen[4], t73, t63, t53, t43, carry[3]);
AN5 A3A(carry_in, tr[7], tr[6], tr[5], tr[4], t73);
AN4 A3B(gen[7], tr[6], tr[5], tr[4], t63);
AN3 A3C(gen[6], tr[5], tr[4], t53);
AN2 A3D(gen[5], tr[4], t43);
OR2 CY2A(t42, t32, t4232);
OR5 CY2(gen[3], t72, t62, t52, t4232, carry[2]);
AN2 A2AA(tr[4], tr[3], tr43);
AN5 A2A(carry_in, tr[7], tr[6], tr[5], tr43, t72);
AN4 A2B(gen[7], tr[6], tr[5], tr43, t62);
AN3 A2C(gen[6], tr[5], tr43, t52);
AN2 A2D(gen[5], tr43, t42);
AN2 A2E(gen[4], tr[3], t32);
OR3 CY1A(t41, t31, t21, t413121);
OR5 CY1(gen[2], t71, t61, t51, t413121, carry[1]);
AN3 A1AA(tr[4], tr[3], tr[2], tr432);
AN5 A1A(carry_in, tr[7], tr[6], tr[5], tr432, t71);
AN4 A1B(gen[7], tr[6], tr[5], tr432, t61);
AN3 A1C(gen[6], tr[5], tr432, t51);
AN2 A1D(gen[5], tr432, t41);
AN3 A1E(gen[4], tr[3], tr[2], t31);
AN2 A1F(gen[3], tr[2], t21);
OR4 CY0A(t40, t30, t20, t10, t40302010);
OR5 CY0(gen[1], t70, t60, t50, t40302010, carry[0]);
AN4 A0AA(tr[4], tr[3], tr[2], tr[1], tr4321);
AN5 A0A(carry_in, tr[7], tr[6], tr[5], tr4321, t70);
AN4 A0B(gen[7], tr[6], tr[5], tr4321, t60);
AN3 A0C(gen[6], tr[5], tr4321, t50);
AN2 A0D(gen[5], tr4321, t40);
AN4 A0E(gen[4], tr[3], tr[2], tr[1], t30);
AN3 A0F(gen[3], tr[2], tr[1], t20);
AN2 A0G(gen[2], tr[1], t10);
OR4 GCYA(t4g, t3g, t2g, t1g, t4321g);
OR5 GCY(gen[0], t7g, t6g, t5g, t4321g, ggen);
AN5 AgA(gen[7], tr[6], tr[5], tr4321, tr[0], t7g);
AN4 AgB(gen[6], tr[5], tr4321, tr[0], t6g);
AN3 AgC(gen[5], tr4321, tr[0], t5g);
AN5 AgD(gen[4], tr[3], tr[2], tr[1], tr[0], t4g);
AN4 AgE(gen[3], tr[2], tr[1], tr[0], t3g);
AN3 AgF(gen[2], tr[1], tr[0], t2g);
AN2 AgG(gen[1], tr[0], t1g);
AN5 GTR(tr[7], tr[6], tr[5], tr4321, tr[0], gtran);

endmodule

// End of DAS Multipier circuit
