module	OR3(a, b, c, z);

input	a, b, c;
output	z;

or #1 g1(z, a, b, c);

endmodule
