module	AN3(a, b, c, z);

input	a, b, c;
output	z;

and #1 g1(z, a, b, c);

endmodule
