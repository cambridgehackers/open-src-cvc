// C880.blif
module foobar(i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1);
input a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1;
output i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2;
not(i2, h1);
and(j2, c1, g1);
and(k2, c1, e1);
and(l2, c1, d1);
or(m2, v0, u0);
not(t_0, v0);
not(t_1, u0);
or(n2, t_0, t_1);
or(o2, t0, s0);
not(t_2, t0);
not(t_3, s0);
or(p2, t_2, t_3);
or(q2, r0, q0);
not(t_4, r0);
not(t_5, q0);
or(r2, t_4, t_5);
or(s2, p0, o0);
not(t_6, p0);
not(t_7, o0);
or(t2, t_6, t_7);
and(u2, l0, h0);
and(v2, x0, d0);
or(w2, e0, d0);
not(t_8, e0);
not(t_9, d0);
or(x2, t_8, t_9);
and(y2, x0, c0);
and(z2, x0, b0);
or(a3, c0, b0);
not(t_10, c0);
not(t_11, b0);
or(b3, t_10, t_11);
and(c3, x0, a0);
and(d3, x0, z);
or(e3, a0, z);
not(t_12, a0);
not(t_13, z);
or(f3, t_12, t_13);
and(g3, x0, y);
and(h3, x0, x);
or(i3, y, x);
not(t_14, y);
not(t_15, x);
or(j3, t_14, t_15);
or(k3, u, t);
and(l1, r, s);
not(t_16, n0);
not(t_17, k);
or(m3, t_16, t_17);
and(n3, k, p, q);
not(t_18, o);
not(t_19, l);
not(t_20, k);
or(o3, t_18, t_19, t_20);
and(p3, i, h0);
and(q3, k, p, h);
not(t_21, m);
not(t_22, l);
not(t_23, h);
not(t_24, k);
or(r3, t_21, t_22, t_23, t_24);
and(s3, k, g, h);
and(t3, k, g, q);
and(k1, f, g, h);
and(j1, f, g, q);
and(i1, f, p, h);
and(x3, f, p, q);
not(t_25, l);
not(t_26, f);
or(y3, t_25, t_26);
and(z3, f, g, h);
and(a4, d, h);
not(t_27, d);
not(t_28, h);
and(b4, t_27, t_28);
and(c4, d, h0);
and(d4, b, h0);
not(t_29, j);
not(t_30, c);
not(t_31, b);
not(t_32, a);
or(e4, t_29, t_30, t_31, t_32);
not(t_33, d);
not(t_34, i);
not(t_35, b);
not(t_36, a);
or(f4, t_33, t_34, t_35, t_36);
and(g4, a, e, i);
not(t_37, d);
not(t_38, c);
not(t_39, e);
not(t_40, a);
or(h4, t_37, t_38, t_39, t_40);
not(t_41, d);
not(t_42, c);
not(t_43, b);
not(t_44, a);
or(i4, t_41, t_42, t_43, t_44);
not(j4, i2);
not(t_45, m2);
not(t_46, n2);
or(k4, t_45, t_46);
not(t_47, o2);
not(t_48, p2);
or(l4, t_47, t_48);
not(t_49, q2);
not(t_50, r2);
or(m4, t_49, t_50);
not(t_51, s2);
not(t_52, t2);
or(n4, t_51, t_52);
not(t_53, w2);
not(t_54, x2);
or(o4, t_53, t_54);
not(t_55, a3);
not(t_56, b3);
or(p4, t_55, t_56);
not(t_57, e3);
not(t_58, f3);
or(q4, t_57, t_58);
not(t_59, i3);
not(t_60, j3);
or(r4, t_59, t_60);
and(r1, w, k3);
not(t_61, k3);
not(t_62, v);
or(t4, t_61, t_62);
not(o1, n3);
or(v4, o3, e4);
not(w4, q3);
not(t_63, e4);
not(t_64, r3);
and(x4, t_63, t_64);
not(q1, s3);
not(p1, t3);
or(a5, y3, e4);
not(b5, z3);
or(n1, z3, h4);
not(t_65, b4);
not(t_66, a4);
and(d5, t_65, t_66);
not(e5, f4);
not(f5, g4);
not(g5, g4);
not(m1, i4);
and(i5, x0, j4);
not(j5, k4);
and(k5, l4, k4);
not(l5, l4);
not(m5, m4);
and(n5, n4, m4);
not(o5, n4);
not(p5, o4);
and(q5, p4, o4);
not(r5, p4);
not(s5, q4);
and(t5, r4, q4);
not(u5, r4);
not(w1, t4);
and(w5, x4, n);
not(v1, v4);
not(t_67, w4);
not(t_68, e5);
or(y5, t_67, t_68);
not(u1, a5);
not(a6, f5);
not(t1, g5);
or(s1, b5, h4);
and(d6, l5, j5);
and(e6, o5, m5);
and(f6, r5, p5);
and(g6, u5, s5);
not(h6, w5);
not(t_69, a6);
not(t_70, n0);
not(t_71, k);
not(t_72, d5);
or(i6, t_69, t_70, t_71, t_72);
not(t_73, j);
not(t_74, x3);
not(t_75, a6);
or(j6, t_73, t_74, t_75);
and(k6, m3, a6, j);
not(t_76, d);
not(t_77, m3);
not(t_78, a6);
or(l6, t_76, t_77, t_78);
and(m6, a6, d, x3);
or(n6, j6, j4);
or(o6, j6, j4);
or(p6, j6, j4);
or(q6, j6, j4);
and(r6, i2, m6);
and(s6, i2, m6);
and(t6, i2, m6);
and(u6, i2, m6);
not(t_79, k5);
not(t_80, d6);
and(v6, t_79, t_80);
not(t_81, n5);
not(t_82, e6);
and(w6, t_81, t_82);
and(x6, m0, k6);
and(y6, k0, k6);
and(z6, j0, k6);
and(a7, i0, k6);
not(t_83, q5);
not(t_84, f6);
and(b7, t_83, t_84);
not(t_85, t5);
not(t_86, g6);
and(c7, t_85, t_86);
not(d7, h6);
not(t_87, y5);
not(t_88, i6);
or(e7, t_87, t_88);
not(t_89, a);
not(t_90, l6);
or(f7, t_89, t_90);
not(t_91, a7);
not(t_92, r6);
and(g7, t_91, t_92);
not(t_93, z6);
not(t_94, s6);
and(h7, t_93, t_94);
not(t_95, y6);
not(t_96, t6);
and(i7, t_95, t_96);
not(t_97, x6);
not(t_98, u6);
and(j7, t_97, t_98);
or(k7, w0, v6);
not(t_99, w0);
not(t_100, v6);
or(l7, t_99, t_100);
not(t_101, v0);
not(t_102, d7);
or(m7, t_101, t_102);
not(t_103, u0);
not(t_104, d7);
or(n7, t_103, t_104);
not(t_105, t0);
not(t_106, d7);
or(o7, t_105, t_106);
and(p7, d7, s0);
and(q7, d7, r0);
and(r7, d7, q0);
and(s7, d7, p0);
and(t7, d7, o0);
and(u7, m0, f7);
and(v7, k0, f7);
and(w7, j0, f7);
and(x7, i0, f7);
or(y7, g0, b7);
not(t_107, g0);
not(t_108, b7);
or(z7, t_107, t_108);
or(a8, w6, f0);
not(t_109, w6);
not(t_110, f0);
or(b8, t_109, t_110);
or(c8, c7, f0);
not(t_111, c7);
not(t_112, f0);
or(d8, t_111, t_112);
and(e8, e0, e7);
and(f8, d0, e7);
and(g8, c0, e7);
and(h8, b0, e7);
and(i8, a0, e7);
and(j8, z, e7);
and(k8, y, e7);
and(l8, x, e7);
not(t_113, k7);
not(t_114, l7);
or(m8, t_113, t_114);
not(t_115, u7);
not(t_116, e8);
and(n8, t_115, t_116);
not(t_117, v7);
not(t_118, f8);
and(o8, t_117, t_118);
not(t_119, w7);
not(t_120, g8);
and(p8, t_119, t_120);
not(t_121, x7);
not(t_122, h8);
and(q8, t_121, t_122);
not(t_123, u2);
not(t_124, i8);
and(r8, t_123, t_124);
not(t_125, y7);
not(t_126, z7);
or(s8, t_125, t_126);
not(t_127, a8);
not(t_128, b8);
or(t8, t_127, t_128);
not(t_129, c8);
not(t_130, d8);
or(u8, t_129, t_130);
not(t_131, p3);
not(t_132, k8);
and(v8, t_131, t_132);
not(t_133, c4);
not(t_134, j8);
and(w8, t_133, t_134);
not(t_135, d4);
not(t_136, l8);
and(x8, t_135, t_136);
not(t_137, q8);
not(t_138, n6);
or(y8, t_137, t_138);
not(t_139, p8);
not(t_140, o6);
or(z8, t_139, t_140);
not(t_141, o8);
not(t_142, p6);
or(a9, t_141, t_142);
not(t_143, n8);
not(t_144, q6);
or(b9, t_143, t_144);
not(t_145, g7);
not(t_146, x8);
or(c9, t_145, t_146);
not(t_147, h7);
not(t_148, v8);
or(d9, t_147, t_148);
not(t_149, i7);
not(t_150, w8);
or(e9, t_149, t_150);
not(t_151, j7);
not(t_152, r8);
or(f9, t_151, t_152);
not(g9, m8);
and(h9, t8, m8);
not(i9, s8);
and(j9, u8, s8);
not(k9, t8);
not(l9, u8);
and(m9, b1, b9);
and(n9, b1, a9);
and(o9, b1, z8);
and(p9, b1, y8);
and(q9, b1, f9);
and(r9, b1, e9);
and(s9, b1, d9);
and(t9, b1, c9);
and(u9, k9, g9);
or(v9, v0, b9);
not(t_153, v0);
not(t_154, b9);
or(w9, t_153, t_154);
or(x9, u0, a9);
not(t_155, u0);
not(t_156, a9);
or(y9, t_155, t_156);
or(z9, t0, z8);
not(t_157, t0);
not(t_158, z8);
or(a10, t_157, t_158);
or(b10, s0, y8);
not(t_159, s0);
not(t_160, y8);
or(c10, t_159, t_160);
or(d10, r0, f9);
not(t_161, r0);
not(t_162, f9);
or(e10, t_161, t_162);
or(f10, q0, e9);
not(t_163, q0);
not(t_164, e9);
or(g10, t_163, t_164);
or(h10, p0, d9);
not(t_165, p0);
not(t_166, d9);
or(i10, t_165, t_166);
or(j10, o0, c9);
not(t_167, o0);
not(t_168, c9);
or(k10, t_167, t_168);
and(l10, l9, i9);
not(t_169, f1);
not(t_170, v9);
not(t_171, x9);
not(t_172, z9);
or(m10, t_169, t_170, t_171, t_172);
not(t_173, f1);
not(t_174, v9);
not(t_175, x9);
or(n10, t_173, t_174, t_175);
not(t_176, f1);
not(t_177, v9);
or(o10, t_176, t_177);
not(t_178, j2);
not(t_179, m9);
and(p10, t_178, t_179);
not(t_180, k2);
not(t_181, n9);
and(q10, t_180, t_181);
not(t_182, l2);
not(t_183, o9);
and(r10, t_182, t_183);
not(t_184, h9);
not(t_185, u9);
and(y1, t_184, t_185);
and(t10, v9, w9);
not(u10, w9);
and(v10, x9, y9);
not(w10, y9);
and(x10, z9, a10);
not(y10, a10);
and(z10, b10, c10);
not(a11, c10);
not(t_186, p9);
not(t_187, p7);
and(b11, t_186, t_187);
and(c11, d10, e10);
not(d11, e10);
not(t_188, q9);
not(t_189, q7);
and(e11, t_188, t_189);
and(f11, f10, g10);
not(g11, g10);
not(t_190, r9);
not(t_191, r7);
and(h11, t_190, t_191);
and(i11, h10, i10);
not(j11, i10);
not(t_192, s9);
not(t_193, s7);
and(k11, t_192, t_193);
and(l11, j10, k10);
not(m11, k10);
not(t_194, t9);
not(t_195, t7);
and(n11, t_194, t_195);
not(t_196, j9);
not(t_197, l10);
and(x1, t_196, t_197);
and(p11, t10, f1);
not(t_198, t10);
not(t_199, f1);
and(q11, t_198, t_199);
and(r11, a1, u10);
and(s11, a1, w10);
and(t11, a1, y10);
and(u11, a1, a11);
and(v11, a1, d11);
and(w11, a1, g11);
and(x11, a1, j11);
and(y11, a1, m11);
and(z11, z0, t10);
and(a12, z0, v10);
and(b12, z0, x10);
and(c12, z0, z10);
and(d12, z0, c11);
and(e12, z0, f11);
and(f12, z0, i11);
and(g12, z0, l11);
not(h12, u10);
not(t_200, u10);
not(t_201, x9);
or(i12, t_200, t_201);
not(t_202, u10);
not(t_203, x9);
not(t_204, z9);
or(j12, t_202, t_203, t_204);
not(k12, w10);
not(t_205, w10);
not(t_206, z9);
or(l12, t_205, t_206);
not(m12, y10);
not(n12, a11);
not(o12, d11);
not(t_207, d11);
not(t_208, f10);
or(p12, t_207, t_208);
not(t_209, d11);
not(t_210, f10);
not(t_211, h10);
or(q12, t_209, t_210, t_211);
not(r12, g11);
not(t_212, g11);
not(t_213, h10);
or(s12, t_212, t_213);
not(t12, j11);
not(u12, m11);
not(t_214, q11);
not(t_215, p11);
and(v12, t_214, t_215);
not(t_216, m10);
not(t_217, j12);
not(t_218, l12);
not(t_219, m12);
or(w12, t_216, t_217, t_218, t_219);
not(t_220, n10);
not(t_221, i12);
not(t_222, k12);
or(x12, t_220, t_221, t_222);
not(t_223, o10);
not(t_224, h12);
or(y12, t_223, t_224);
not(t_225, z11);
not(t_226, r11);
and(z12, t_225, t_226);
not(t_227, a12);
not(t_228, s11);
and(a13, t_227, t_228);
not(t_229, b12);
not(t_230, t11);
and(b13, t_229, t_230);
not(t_231, c12);
not(t_232, u11);
and(c13, t_231, t_232);
not(t_233, d12);
not(t_234, v11);
and(d13, t_233, t_234);
not(t_235, e12);
not(t_236, w11);
and(e13, t_235, t_236);
not(t_237, f12);
not(t_238, x11);
and(f13, t_237, t_238);
not(t_239, g12);
not(t_240, y11);
and(g13, t_239, t_240);
and(h13, y0, v12);
not(t_241, v10);
not(t_242, y12);
and(i13, t_241, t_242);
and(j13, v10, y12);
not(t_243, x10);
not(t_244, x12);
and(k13, t_243, t_244);
and(l13, x10, x12);
not(t_245, z10);
not(t_246, w12);
and(m13, t_245, t_246);
and(n13, z10, w12);
not(t_247, w12);
not(t_248, b10);
or(o13, t_247, t_248);
not(t_249, i13);
not(t_250, j13);
and(p13, t_249, t_250);
not(t_251, k13);
not(t_252, l13);
and(q13, t_251, t_252);
not(t_253, m13);
not(t_254, n13);
and(r13, t_253, t_254);
not(t_255, n12);
not(t_256, o13);
or(s13, t_255, t_256);
not(t_257, v2);
not(t_258, h13);
and(t13, t_257, t_258);
and(u13, y0, p13);
and(v13, y0, q13);
and(w13, y0, r13);
not(t_259, m7);
not(t_260, p10);
not(t_261, z12);
not(t_262, t13);
or(x13, t_259, t_260, t_261, t_262);
not(t_263, c11);
not(t_264, s13);
and(y13, t_263, t_264);
and(z13, c11, s13);
not(t_265, s13);
not(t_266, d10);
or(a14, t_265, t_266);
not(t_267, s13);
not(t_268, d10);
not(t_269, f10);
or(b14, t_267, t_268, t_269);
not(t_270, s13);
not(t_271, d10);
not(t_272, f10);
not(t_273, h10);
or(c14, t_270, t_271, t_272, t_273);
not(d14, x13);
not(t_274, y13);
not(t_275, z13);
and(e14, t_274, t_275);
not(t_276, a14);
not(t_277, o12);
or(f14, t_276, t_277);
not(t_278, b14);
not(t_279, p12);
not(t_280, r12);
or(g14, t_278, t_279, t_280);
not(t_281, c14);
not(t_282, q12);
not(t_283, s12);
not(t_284, t12);
or(h14, t_281, t_282, t_283, t_284);
not(t_285, y2);
not(t_286, u13);
and(i14, t_285, t_286);
not(t_287, z2);
not(t_288, v13);
and(j14, t_287, t_288);
not(t_289, c3);
not(t_290, w13);
and(k14, t_289, t_290);
and(l14, y0, e14);
not(z1, d14);
not(t_291, n7);
not(t_292, q10);
not(t_293, a13);
not(t_294, i14);
or(n14, t_291, t_292, t_293, t_294);
not(t_295, o7);
not(t_296, r10);
not(t_297, b13);
not(t_298, j14);
or(o14, t_295, t_296, t_297, t_298);
not(t_299, b11);
not(t_300, c13);
not(t_301, k14);
or(p14, t_299, t_300, t_301);
not(t_302, f11);
not(t_303, f14);
and(q14, t_302, t_303);
and(r14, f11, f14);
not(t_304, i11);
not(t_305, g14);
and(s14, t_304, t_305);
and(t14, i11, g14);
not(t_306, l11);
not(t_307, h14);
and(u14, t_306, t_307);
and(v14, l11, h14);
not(t_308, j10);
not(t_309, h14);
or(w14, t_308, t_309);
not(x14, n14);
not(y14, o14);
not(z14, p14);
not(t_310, q14);
not(t_311, r14);
and(a15, t_310, t_311);
not(t_312, s14);
not(t_313, t14);
and(b15, t_312, t_313);
not(t_314, u14);
not(t_315, v14);
and(c15, t_314, t_315);
and(d15, u12, w14);
not(t_316, d3);
not(t_317, l14);
and(e15, t_316, t_317);
and(f15, y0, a15);
and(g15, y0, b15);
and(h15, y0, c15);
not(c2, x14);
not(b2, y14);
not(a2, z14);
not(t_318, e11);
not(t_319, d13);
not(t_320, e15);
or(l15, t_318, t_319, t_320);
not(d2, d15);
not(t_321, i5);
not(t_322, h15);
and(n15, t_321, t_322);
not(o15, l15);
not(t_323, g3);
not(t_324, f15);
and(p15, t_323, t_324);
not(t_325, h3);
not(t_326, g15);
and(q15, t_325, t_326);
not(e2, o15);
not(t_327, h11);
not(t_328, e13);
not(t_329, p15);
or(s15, t_327, t_328, t_329);
not(t_330, k11);
not(t_331, f13);
not(t_332, q15);
or(t15, t_330, t_331, t_332);
not(t_333, n11);
not(t_334, g13);
not(t_335, n15);
or(u15, t_333, t_334, t_335);
not(v15, s15);
not(w15, t15);
not(x15, u15);
not(h2, v15);
not(g2, w15);
not(f2, x15);
endmodule
module top;
	parameter in_width = 60,
		// patterns = 5000,
		patterns = 8,
		step = 1;
	reg [1:in_width] in_mem[1:patterns];
	integer index;

	wire i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
		i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,
		i50,i51,i52,i53,i54,i55,i56,i57,i58,i59;

	assign {i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
		i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,
		i50,i51,i52,i53,i54,i55,i56,i57,i58,i59} = 
		$getpattern(in_mem[index]);

	initial $monitor($time,,o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,
		o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
		o20,o21,o22,o23,o24,o25);
	initial
		begin
			$readmemb("patt.mem", in_mem);
			for(index = 1; index <= patterns; index = index + 1)
				#step;
		end

	foobar cct(o0,o1,o2,o3,o4,o5,o6,o7,o8,o9,
		o10,o11,o12,o13,o14,o15,o16,o17,o18,o19,
		o20,o21,o22,o23,o24,o25,i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,
		i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
		i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
		i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
		i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,
		i50,i51,i52,i53,i54,i55,i56,i57,i58,i59);
endmodule
