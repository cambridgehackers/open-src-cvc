module	AN4(a, b, c, d, z);

input	a, b, c, d;
output	z;

and #1 g1(z, a, b, c, d);

endmodule
